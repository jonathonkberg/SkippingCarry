* SPICE NETLIST
***************************************

.SUBCKT i
** N=13 EP=0 IP=0 FDC=0
* PORT VDD VDD -23500 1500 METAL2
* PORT IN2 IN2 -21000 30000 METAL1
* PORT IN2 IN2 151000 58000 METAL1
* PORT IN4 IN4 -21000 44000 METAL1
* PORT IN4 IN4 151000 30000 METAL1
* PORT IN3 IN3 -21000 58000 METAL1
* PORT IN3 IN3 151000 44000 METAL1
* PORT IN1 IN1 -21000 72000 METAL1
* PORT IN1 IN1 151000 72000 METAL1
* PORT OUTN OUTN 37000 -33000 METAL1
* PORT OUT OUT 79000 -33000 METAL1
* PORT GND GND 151000 10000 METAL1
*.SEEDPROM
.ENDS
***************************************
.SUBCKT full_adder GND COUTN COUT VDD BN A CN C P B AN
** N=32 EP=11 IP=52 FDC=44
* PORT SUM <UNATTACHED> -176951 131998 <UNATTACHED>
* PORT COUTN <UNATTACHED> 533349 216244 <UNATTACHED>
* PORT GND GND 715667 191032 METAL1
* PORT COUTN GND 718086 191561 METAL1
* PORT COUTN COUTN 412148 113156 METAL1
* PORT COUT COUT 454492 113156 METAL1
* PORT VDD VDD -176088 182434 METAL2
* PORT BN BN 715652 210954 METAL1
* PORT A A 715693 252942 METAL1
* PORT CN CN 412507 316865 METAL1
* PORT C C 454647 298940 METAL1
* PORT P P 640803 131375 METAL1
* PORT B B 715687 224942 METAL1
* PORT AN AN 715707 238986 METAL1
M0 GND 8 10 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=134209 $Y=180008 $D=1
M1 GND 5 8 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=137209 $Y=224008 $D=1
M2 27 6 GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=137209 $Y=238008 $D=1
M3 8 BN 27 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=137209 $Y=252008 $D=1
M4 GND 5 A GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=281565 $Y=197014 $D=1
M5 5 6 GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=292565 $Y=238014 $D=1
M6 GND BN 5 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=292565 $Y=252014 $D=1
M7 GND 18 19 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=-63099 $Y=168994 $D=1
M8 GND COUTN COUT GND N L=2.0124e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=465049 $Y=183000 $D=1
M9 GND 23 P GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=654684 $Y=168964 $D=1
M10 25 P 18 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=-40099 $Y=209994 $D=1
M11 28 6 COUTN GND N L=2.0124e-07 W=5.4e-07 AD=5.7173e-13 AS=4.374e-13 $X=488049 $Y=224000 $D=1
M12 30 BN 23 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=677684 $Y=209964 $D=1
M13 GND 10 25 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=-40099 $Y=223994 $D=1
M14 GND BN 28 GND N L=2.0124e-07 W=5.4e-07 AD=5.7173e-13 AS=5.7173e-13 $X=488049 $Y=238000 $D=1
M15 GND B 30 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=677684 $Y=223964 $D=1
M16 26 C GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=-40099 $Y=237994 $D=1
M17 29 A GND GND N L=2.0124e-07 W=5.4e-07 AD=5.7173e-13 AS=5.7173e-13 $X=488049 $Y=252000 $D=1
M18 31 AN GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=677684 $Y=237964 $D=1
M19 18 CN 26 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=-40099 $Y=251994 $D=1
M20 COUTN 20 29 GND N L=2.0124e-07 W=5.4e-07 AD=4.374e-13 AS=5.7173e-13 $X=488049 $Y=266000 $D=1
M21 23 A 31 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=677684 $Y=251964 $D=1
M22 9 5 8 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=78209 $Y=224008 $D=0
M23 VDD 6 9 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=78209 $Y=238008 $D=0
M24 9 BN VDD VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=78209 $Y=252008 $D=0
M25 VDD 8 10 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=93209 $Y=180008 $D=0
M26 32 6 VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=231565 $Y=238014 $D=0
M27 5 BN 32 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=231565 $Y=252014 $D=0
M28 VDD 5 A VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=247565 $Y=197014 $D=0
M29 VDD 18 19 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-104099 $Y=168994 $D=0
M30 VDD COUTN COUT VDD P L=2.0124e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=424049 $Y=183000 $D=0
M31 VDD 23 P VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=613684 $Y=168964 $D=0
M32 17 C VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=-120099 $Y=209994 $D=0
M33 21 A VDD VDD P L=2.0124e-07 W=2.88e-06 AD=3.04923e-12 AS=2.3328e-12 $X=408049 $Y=224000 $D=0
M34 22 AN VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=597684 $Y=209964 $D=0
M35 18 P 17 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=-120099 $Y=223994 $D=0
M36 COUTN 6 21 VDD P L=2.0124e-07 W=2.88e-06 AD=3.04923e-12 AS=3.04923e-12 $X=408049 $Y=238000 $D=0
M37 23 BN 22 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=597684 $Y=223964 $D=0
M38 17 10 18 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=-120099 $Y=237994 $D=0
M39 21 BN COUTN VDD P L=2.0124e-07 W=2.88e-06 AD=3.04923e-12 AS=3.04923e-12 $X=408049 $Y=252000 $D=0
M40 22 B 23 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=597684 $Y=237964 $D=0
M41 VDD CN 17 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=-120099 $Y=251994 $D=0
M42 VDD 20 21 VDD P L=2.0124e-07 W=2.88e-06 AD=2.3328e-12 AS=3.04923e-12 $X=408049 $Y=266000 $D=0
M43 VDD A 22 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=597684 $Y=251964 $D=0
.ENDS
***************************************
