* Inverter Pre Layout Sub-circuit
* Dec 2022

.include /afs/cad/u/j/k/jk526/ece658/final_project/pre_sim/subckts/inverter_180nm.sp

.subckt sub_ii INI IN2 IN3 IN4 IN5 IN6 OUTN OUT vdd gnd



x1 OUTN OUT vdd gnd INV

.ends
