* File: thirty_two_bit_adder.pex.netlist
* Created: Mon Dec 19 17:36:08 2022
* Program "Calibre xRC"
* Version "v2012.2_36.25"
* 
.include "thirty_two_bit_adder.pex.netlist.pex"
.subckt THIRTY_TWO_BIT_ADDER  VDD COUT31N C0N GND SUM30 SUM26 SUM22 SUM29 SUM25
+ SUM21 SUM28 SUM24 SUM20 SUM31 SUM27 SUM23 SUM14 SUM10 SUM18 SUM6 SUM13 SUM9
+ SUM17 SUM5 SUM12 SUM8 SUM16 SUM4 SUM15 SUM11 SUM19 SUM7 SUM2 SUM1 SUM0 SUM3
+ COUT31 C0 A30N B30 B30N A30 A26N B26 B26N A26 A22N B22 B22N A22 A29N B29 B29N
+ A29 A25N B25 B25N A25 A21N B21 B21N A21 A28N B28 B28N A28 A24N B24 B24N A24
+ A20N B20 B20N A20 A31N B31 B31N A31 A27N B27 B27N A27 A23N B23 B23N A23 A14N
+ B14 B14N A14 A10N B10 B10N A10 A18N B18 B18N A18 A6N B6 B6N A6 A13N B13 B13N
+ A13 A9N B9 B9N A9 A17N B17 B17N A17 A5N B5 B5N A5 A12N B12 B12N A12 A8N B8 B8N
+ A8 A16N B16 B16N A16 A4N B4 B4N A4 A15N B15 B15N A15 A11N B11 B11N A11 A19N
+ B19 B19N A19 A7N B7 B7N A7 A2N B2 B2N A2 A1N B1 B1N A1 A0N B0 B0N A0 A3N B3
+ B3N A3
* 
* A3	A3
* B3N	B3N
* B3	B3
* A3N	A3N
* A0	A0
* B0N	B0N
* B0	B0
* A0N	A0N
* A1	A1
* B1N	B1N
* B1	B1
* A1N	A1N
* A2	A2
* B2N	B2N
* B2	B2
* A2N	A2N
* A7	A7
* B7N	B7N
* B7	B7
* A7N	A7N
* A19	A19
* B19N	B19N
* B19	B19
* A19N	A19N
* A11	A11
* B11N	B11N
* B11	B11
* A11N	A11N
* A15	A15
* B15N	B15N
* B15	B15
* A15N	A15N
* A4	A4
* B4N	B4N
* B4	B4
* A4N	A4N
* A16	A16
* B16N	B16N
* B16	B16
* A16N	A16N
* A8	A8
* B8N	B8N
* B8	B8
* A8N	A8N
* A12	A12
* B12N	B12N
* B12	B12
* A12N	A12N
* A5	A5
* B5N	B5N
* B5	B5
* A5N	A5N
* A17	A17
* B17N	B17N
* B17	B17
* A17N	A17N
* A9	A9
* B9N	B9N
* B9	B9
* A9N	A9N
* A13	A13
* B13N	B13N
* B13	B13
* A13N	A13N
* A6	A6
* B6N	B6N
* B6	B6
* A6N	A6N
* A18	A18
* B18N	B18N
* B18	B18
* A18N	A18N
* A10	A10
* B10N	B10N
* B10	B10
* A10N	A10N
* A14	A14
* B14N	B14N
* B14	B14
* A14N	A14N
* A23	A23
* B23N	B23N
* B23	B23
* A23N	A23N
* A27	A27
* B27N	B27N
* B27	B27
* A27N	A27N
* A31	A31
* B31N	B31N
* B31	B31
* A31N	A31N
* A20	A20
* B20N	B20N
* B20	B20
* A20N	A20N
* A24	A24
* B24N	B24N
* B24	B24
* A24N	A24N
* A28	A28
* B28N	B28N
* B28	B28
* A28N	A28N
* A21	A21
* B21N	B21N
* B21	B21
* A21N	A21N
* A25	A25
* B25N	B25N
* B25	B25
* A25N	A25N
* A29	A29
* B29N	B29N
* B29	B29
* A29N	A29N
* A22	A22
* B22N	B22N
* B22	B22
* A22N	A22N
* A26	A26
* B26N	B26N
* B26	B26
* A26N	A26N
* A30	A30
* B30N	B30N
* B30	B30
* A30N	A30N
* C0	C0
* COUT31	COUT31
* SUM3	SUM3
* SUM0	SUM0
* SUM1	SUM1
* SUM2	SUM2
* SUM7	SUM7
* SUM19	SUM19
* SUM11	SUM11
* SUM15	SUM15
* SUM4	SUM4
* SUM16	SUM16
* SUM8	SUM8
* SUM12	SUM12
* SUM5	SUM5
* SUM17	SUM17
* SUM9	SUM9
* SUM13	SUM13
* SUM6	SUM6
* SUM18	SUM18
* SUM10	SUM10
* SUM14	SUM14
* SUM23	SUM23
* SUM27	SUM27
* SUM31	SUM31
* SUM20	SUM20
* SUM24	SUM24
* SUM28	SUM28
* SUM21	SUM21
* SUM25	SUM25
* SUM29	SUM29
* SUM22	SUM22
* SUM26	SUM26
* SUM30	SUM30
* GND	GND
* C0N	C0N
* COUT31N	COUT31N
* VDD	VDD
mX0/M0 N_GND_X0/M0_d N_X0/39_X0/M0_g N_X0/40_X0/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/M1 N_X0/41_X0/M1_d N_X0/32_X0/M1_g N_GND_X0/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX0/M2 N_X0/42_X0/M2_d N_X0/31_X0/M2_g N_X0/41_X0/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX0/M3 N_X0/43_X0/M3_d N_X0/30_X0/M3_g N_X0/42_X0/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX0/M4 N_X0/39_X0/M4_d N_X0/35_X0/M4_g N_X0/43_X0/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX0/M5 N_VDD_X0/M5_d N_X0/39_X0/M5_g N_X0/40_X0/M5_s N_VDD_X0/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/M6 N_X0/39_X0/M6_d N_X0/32_X0/M6_g N_VDD_X0/M6_s N_VDD_X0/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX0/M7 N_VDD_X0/M7_d N_X0/31_X0/M7_g N_X0/39_X0/M7_s N_VDD_X0/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX0/M8 N_X0/39_X0/M8_d N_X0/30_X0/M8_g N_VDD_X0/M8_s N_VDD_X0/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX0/M9 N_VDD_X0/M9_d N_X0/35_X0/M9_g N_X0/39_X0/M9_s N_VDD_X0/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX0/X10/M0 N_GND_X0/X10/M0_d N_COUT31N_X0/X10/M0_g N_COUT31_X0/X10/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X10/M1 N_X0/X10/10_X0/X10/M1_d N_45_X0/X10/M1_g N_COUT31N_X0/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X10/M2 N_GND_X0/X10/M2_d N_X0/40_X0/X10/M2_g N_X0/X10/10_X0/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X10/M3 N_X0/X10/11_X0/X10/M3_d N_X0/39_X0/X10/M3_g N_GND_X0/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X10/M4 N_COUT31N_X0/X10/M4_d N_X0/34_X0/X10/M4_g N_X0/X10/11_X0/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X10/M5 N_X0/X10/9_X0/X10/M5_d N_X0/39_X0/X10/M5_g N_VDD_X0/X10/M5_s
+ N_VDD_X0/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX0/X10/M6 N_COUT31N_X0/X10/M6_d N_45_X0/X10/M6_g N_X0/X10/9_X0/X10/M6_s
+ N_VDD_X0/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X10/M7 N_X0/X10/9_X0/X10/M7_d N_X0/40_X0/X10/M7_g N_COUT31N_X0/X10/M7_s
+ N_VDD_X0/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X10/M8 N_VDD_X0/X10/M8_d N_X0/34_X0/X10/M8_g N_X0/X10/9_X0/X10/M8_s
+ N_VDD_X0/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X10/M9 N_VDD_X0/X10/M9_d N_COUT31N_X0/X10/M9_g N_COUT31_X0/X10/M9_s
+ N_VDD_X0/X10/M5_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X11/M0 N_GND_X0/X11/M0_d N_X0/X11/14_X0/X11/M0_g N_X0/X11/16_X0/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X11/M1 N_GND_X0/X11/M1_d N_X0/X11/13_X0/X11/M1_g N_X0/X11/14_X0/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X11/M2 N_X0/X11/20_X0/X11/M2_d N_B30_X0/X11/M2_g N_GND_X0/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X11/M3 N_X0/X11/14_X0/X11/M3_d N_A30_X0/X11/M3_g N_X0/X11/20_X0/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X11/M4 N_GND_X0/X11/M4_d N_X0/X11/13_X0/X11/M4_g N_X0/X11/17_X0/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X11/M5 N_X0/X11/13_X0/X11/M5_d N_B30_X0/X11/M5_g N_GND_X0/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X11/M6 N_GND_X0/X11/M6_d N_A30_X0/X11/M6_g N_X0/X11/13_X0/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X11/M7 N_X0/X11/15_X0/X11/M7_d N_X0/X11/13_X0/X11/M7_g
+ N_X0/X11/14_X0/X11/M7_s N_VDD_X0/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX0/X11/M8 N_VDD_X0/X11/M8_d N_B30_X0/X11/M8_g N_X0/X11/15_X0/X11/M8_s
+ N_VDD_X0/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X11/M9 N_X0/X11/15_X0/X11/M9_d N_A30_X0/X11/M9_g N_VDD_X0/X11/M9_s
+ N_VDD_X0/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X11/M10 N_VDD_X0/X11/M10_d N_X0/X11/14_X0/X11/M10_g N_X0/X11/16_X0/X11/M10_s
+ N_VDD_X0/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X11/M11 N_X0/X11/21_X0/X11/M11_d N_B30_X0/X11/M11_g N_VDD_X0/X11/M11_s
+ N_VDD_X0/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX0/X11/M12 N_X0/X11/13_X0/X11/M12_d N_A30_X0/X11/M12_g N_X0/X11/21_X0/X11/M12_s
+ N_VDD_X0/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X11/M13 N_VDD_X0/X11/M13_d N_X0/X11/13_X0/X11/M13_g N_X0/X11/17_X0/X11/M13_s
+ N_VDD_X0/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X11/X14/M0 N_GND_X0/X11/X14/M0_d N_X0/X11/18_X0/X11/X14/M0_g
+ N_SUM30_X0/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X11/X14/M1 N_X0/X11/X14/10_X0/X11/X14/M1_d N_X0/30_X0/X11/X14/M1_g
+ N_X0/X11/18_X0/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X11/X14/M2 N_GND_X0/X11/X14/M2_d N_X0/27_X0/X11/X14/M2_g
+ N_X0/X11/X14/10_X0/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X11/X14/M3 N_X0/X11/X14/11_X0/X11/X14/M3_d N_X0/X11/16_X0/X11/X14/M3_g
+ N_GND_X0/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X11/X14/M4 N_X0/X11/18_X0/X11/X14/M4_d N_X0/36_X0/X11/X14/M4_g
+ N_X0/X11/X14/11_X0/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X11/X14/M5 N_X0/X11/X14/9_X0/X11/X14/M5_d N_X0/X11/16_X0/X11/X14/M5_g
+ N_VDD_X0/X11/X14/M5_s N_VDD_X0/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X11/X14/M6 N_X0/X11/18_X0/X11/X14/M6_d N_X0/30_X0/X11/X14/M6_g
+ N_X0/X11/X14/9_X0/X11/X14/M6_s N_VDD_X0/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X14/M7 N_X0/X11/X14/9_X0/X11/X14/M7_d N_X0/27_X0/X11/X14/M7_g
+ N_X0/X11/18_X0/X11/X14/M7_s N_VDD_X0/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X14/M8 N_VDD_X0/X11/X14/M8_d N_X0/36_X0/X11/X14/M8_g
+ N_X0/X11/X14/9_X0/X11/X14/M8_s N_VDD_X0/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X11/X14/M9 N_VDD_X0/X11/X14/M9_d N_X0/X11/18_X0/X11/X14/M9_g
+ N_SUM30_X0/X11/X14/M9_s N_VDD_X0/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X11/X15/M0 N_GND_X0/X11/X15/M0_d N_X0/29_X0/X11/X15/M0_g
+ N_X0/38_X0/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X11/X15/M1 N_X0/X11/X15/10_X0/X11/X15/M1_d N_X0/X11/17_X0/X11/X15/M1_g
+ N_X0/29_X0/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX0/X11/X15/M2 N_GND_X0/X11/X15/M2_d N_X0/36_X0/X11/X15/M2_g
+ N_X0/X11/X15/10_X0/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X11/X15/M3 N_X0/X11/X15/11_X0/X11/X15/M3_d N_B30_X0/X11/X15/M3_g
+ N_GND_X0/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X11/X15/M4 N_X0/29_X0/X11/X15/M4_d N_A30_X0/X11/X15/M4_g
+ N_X0/X11/X15/11_X0/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X11/X15/M5 N_X0/X11/X15/9_X0/X11/X15/M5_d N_B30_X0/X11/X15/M5_g
+ N_VDD_X0/X11/X15/M5_s N_VDD_X0/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X11/X15/M6 N_X0/29_X0/X11/X15/M6_d N_X0/X11/17_X0/X11/X15/M6_g
+ N_X0/X11/X15/9_X0/X11/X15/M6_s N_VDD_X0/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X15/M7 N_X0/X11/X15/9_X0/X11/X15/M7_d N_X0/36_X0/X11/X15/M7_g
+ N_X0/29_X0/X11/X15/M7_s N_VDD_X0/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X15/M8 N_VDD_X0/X11/X15/M8_d N_A30_X0/X11/X15/M8_g
+ N_X0/X11/X15/9_X0/X11/X15/M8_s N_VDD_X0/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X11/X15/M9 N_VDD_X0/X11/X15/M9_d N_X0/29_X0/X11/X15/M9_g
+ N_X0/38_X0/X11/X15/M9_s N_VDD_X0/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X11/X16/M0 N_GND_X0/X11/X16/M0_d N_X0/X11/19_X0/X11/X16/M0_g
+ N_X0/30_X0/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X11/X16/M1 N_X0/X11/X16/10_X0/X11/X16/M1_d N_A30N_X0/X11/X16/M1_g
+ N_X0/X11/19_X0/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X11/X16/M2 N_GND_X0/X11/X16/M2_d N_B30_X0/X11/X16/M2_g
+ N_X0/X11/X16/10_X0/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X11/X16/M3 N_X0/X11/X16/11_X0/X11/X16/M3_d N_B30N_X0/X11/X16/M3_g
+ N_GND_X0/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X11/X16/M4 N_X0/X11/19_X0/X11/X16/M4_d N_A30_X0/X11/X16/M4_g
+ N_X0/X11/X16/11_X0/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X11/X16/M5 N_X0/X11/X16/9_X0/X11/X16/M5_d N_B30N_X0/X11/X16/M5_g
+ N_VDD_X0/X11/X16/M5_s N_VDD_X0/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X11/X16/M6 N_X0/X11/19_X0/X11/X16/M6_d N_A30N_X0/X11/X16/M6_g
+ N_X0/X11/X16/9_X0/X11/X16/M6_s N_VDD_X0/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X16/M7 N_X0/X11/X16/9_X0/X11/X16/M7_d N_B30_X0/X11/X16/M7_g
+ N_X0/X11/19_X0/X11/X16/M7_s N_VDD_X0/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X11/X16/M8 N_VDD_X0/X11/X16/M8_d N_A30_X0/X11/X16/M8_g
+ N_X0/X11/X16/9_X0/X11/X16/M8_s N_VDD_X0/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X11/X16/M9 N_VDD_X0/X11/X16/M9_d N_X0/X11/19_X0/X11/X16/M9_g
+ N_X0/30_X0/X11/X16/M9_s N_VDD_X0/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X12/M0 N_GND_X0/X12/M0_d N_X0/X12/14_X0/X12/M0_g N_X0/X12/16_X0/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X12/M1 N_GND_X0/X12/M1_d N_X0/X12/13_X0/X12/M1_g N_X0/X12/14_X0/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X12/M2 N_X0/X12/20_X0/X12/M2_d N_B29_X0/X12/M2_g N_GND_X0/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X12/M3 N_X0/X12/14_X0/X12/M3_d N_A29_X0/X12/M3_g N_X0/X12/20_X0/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X12/M4 N_GND_X0/X12/M4_d N_X0/X12/13_X0/X12/M4_g N_X0/X12/17_X0/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X12/M5 N_X0/X12/13_X0/X12/M5_d N_B29_X0/X12/M5_g N_GND_X0/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X12/M6 N_GND_X0/X12/M6_d N_A29_X0/X12/M6_g N_X0/X12/13_X0/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X12/M7 N_X0/X12/15_X0/X12/M7_d N_X0/X12/13_X0/X12/M7_g
+ N_X0/X12/14_X0/X12/M7_s N_VDD_X0/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX0/X12/M8 N_VDD_X0/X12/M8_d N_B29_X0/X12/M8_g N_X0/X12/15_X0/X12/M8_s
+ N_VDD_X0/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X12/M9 N_X0/X12/15_X0/X12/M9_d N_A29_X0/X12/M9_g N_VDD_X0/X12/M9_s
+ N_VDD_X0/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X12/M10 N_VDD_X0/X12/M10_d N_X0/X12/14_X0/X12/M10_g N_X0/X12/16_X0/X12/M10_s
+ N_VDD_X0/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X12/M11 N_X0/X12/21_X0/X12/M11_d N_B29_X0/X12/M11_g N_VDD_X0/X12/M11_s
+ N_VDD_X0/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX0/X12/M12 N_X0/X12/13_X0/X12/M12_d N_A29_X0/X12/M12_g N_X0/X12/21_X0/X12/M12_s
+ N_VDD_X0/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X12/M13 N_VDD_X0/X12/M13_d N_X0/X12/13_X0/X12/M13_g N_X0/X12/17_X0/X12/M13_s
+ N_VDD_X0/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X12/X14/M0 N_GND_X0/X12/X14/M0_d N_X0/X12/18_X0/X12/X14/M0_g
+ N_SUM29_X0/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X12/X14/M1 N_X0/X12/X14/10_X0/X12/X14/M1_d N_X0/31_X0/X12/X14/M1_g
+ N_X0/X12/18_X0/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X12/X14/M2 N_GND_X0/X12/X14/M2_d N_X0/28_X0/X12/X14/M2_g
+ N_X0/X12/X14/10_X0/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X12/X14/M3 N_X0/X12/X14/11_X0/X12/X14/M3_d N_X0/X12/16_X0/X12/X14/M3_g
+ N_GND_X0/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X12/X14/M4 N_X0/X12/18_X0/X12/X14/M4_d N_X0/37_X0/X12/X14/M4_g
+ N_X0/X12/X14/11_X0/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X12/X14/M5 N_X0/X12/X14/9_X0/X12/X14/M5_d N_X0/X12/16_X0/X12/X14/M5_g
+ N_VDD_X0/X12/X14/M5_s N_VDD_X0/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X12/X14/M6 N_X0/X12/18_X0/X12/X14/M6_d N_X0/31_X0/X12/X14/M6_g
+ N_X0/X12/X14/9_X0/X12/X14/M6_s N_VDD_X0/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X14/M7 N_X0/X12/X14/9_X0/X12/X14/M7_d N_X0/28_X0/X12/X14/M7_g
+ N_X0/X12/18_X0/X12/X14/M7_s N_VDD_X0/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X14/M8 N_VDD_X0/X12/X14/M8_d N_X0/37_X0/X12/X14/M8_g
+ N_X0/X12/X14/9_X0/X12/X14/M8_s N_VDD_X0/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X12/X14/M9 N_VDD_X0/X12/X14/M9_d N_X0/X12/18_X0/X12/X14/M9_g
+ N_SUM29_X0/X12/X14/M9_s N_VDD_X0/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X12/X15/M0 N_GND_X0/X12/X15/M0_d N_X0/27_X0/X12/X15/M0_g
+ N_X0/36_X0/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X12/X15/M1 N_X0/X12/X15/10_X0/X12/X15/M1_d N_X0/X12/17_X0/X12/X15/M1_g
+ N_X0/27_X0/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX0/X12/X15/M2 N_GND_X0/X12/X15/M2_d N_X0/37_X0/X12/X15/M2_g
+ N_X0/X12/X15/10_X0/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X12/X15/M3 N_X0/X12/X15/11_X0/X12/X15/M3_d N_B29_X0/X12/X15/M3_g
+ N_GND_X0/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X12/X15/M4 N_X0/27_X0/X12/X15/M4_d N_A29_X0/X12/X15/M4_g
+ N_X0/X12/X15/11_X0/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X12/X15/M5 N_X0/X12/X15/9_X0/X12/X15/M5_d N_B29_X0/X12/X15/M5_g
+ N_VDD_X0/X12/X15/M5_s N_VDD_X0/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X12/X15/M6 N_X0/27_X0/X12/X15/M6_d N_X0/X12/17_X0/X12/X15/M6_g
+ N_X0/X12/X15/9_X0/X12/X15/M6_s N_VDD_X0/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X15/M7 N_X0/X12/X15/9_X0/X12/X15/M7_d N_X0/37_X0/X12/X15/M7_g
+ N_X0/27_X0/X12/X15/M7_s N_VDD_X0/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X15/M8 N_VDD_X0/X12/X15/M8_d N_A29_X0/X12/X15/M8_g
+ N_X0/X12/X15/9_X0/X12/X15/M8_s N_VDD_X0/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X12/X15/M9 N_VDD_X0/X12/X15/M9_d N_X0/27_X0/X12/X15/M9_g
+ N_X0/36_X0/X12/X15/M9_s N_VDD_X0/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X12/X16/M0 N_GND_X0/X12/X16/M0_d N_X0/X12/19_X0/X12/X16/M0_g
+ N_X0/31_X0/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X12/X16/M1 N_X0/X12/X16/10_X0/X12/X16/M1_d N_A29N_X0/X12/X16/M1_g
+ N_X0/X12/19_X0/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X12/X16/M2 N_GND_X0/X12/X16/M2_d N_B29_X0/X12/X16/M2_g
+ N_X0/X12/X16/10_X0/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X12/X16/M3 N_X0/X12/X16/11_X0/X12/X16/M3_d N_B29N_X0/X12/X16/M3_g
+ N_GND_X0/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X12/X16/M4 N_X0/X12/19_X0/X12/X16/M4_d N_A29_X0/X12/X16/M4_g
+ N_X0/X12/X16/11_X0/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X12/X16/M5 N_X0/X12/X16/9_X0/X12/X16/M5_d N_B29N_X0/X12/X16/M5_g
+ N_VDD_X0/X12/X16/M5_s N_VDD_X0/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X12/X16/M6 N_X0/X12/19_X0/X12/X16/M6_d N_A29N_X0/X12/X16/M6_g
+ N_X0/X12/X16/9_X0/X12/X16/M6_s N_VDD_X0/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X16/M7 N_X0/X12/X16/9_X0/X12/X16/M7_d N_B29_X0/X12/X16/M7_g
+ N_X0/X12/19_X0/X12/X16/M7_s N_VDD_X0/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X12/X16/M8 N_VDD_X0/X12/X16/M8_d N_A29_X0/X12/X16/M8_g
+ N_X0/X12/X16/9_X0/X12/X16/M8_s N_VDD_X0/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X12/X16/M9 N_VDD_X0/X12/X16/M9_d N_X0/X12/19_X0/X12/X16/M9_g
+ N_X0/31_X0/X12/X16/M9_s N_VDD_X0/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X13/M0 N_GND_X0/X13/M0_d N_X0/X13/14_X0/X13/M0_g N_X0/X13/16_X0/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X13/M1 N_GND_X0/X13/M1_d N_X0/X13/13_X0/X13/M1_g N_X0/X13/14_X0/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X13/M2 N_X0/X13/20_X0/X13/M2_d N_B28_X0/X13/M2_g N_GND_X0/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X13/M3 N_X0/X13/14_X0/X13/M3_d N_A28_X0/X13/M3_g N_X0/X13/20_X0/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X13/M4 N_GND_X0/X13/M4_d N_X0/X13/13_X0/X13/M4_g N_X0/X13/17_X0/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X13/M5 N_X0/X13/13_X0/X13/M5_d N_B28_X0/X13/M5_g N_GND_X0/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X13/M6 N_GND_X0/X13/M6_d N_A28_X0/X13/M6_g N_X0/X13/13_X0/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X13/M7 N_X0/X13/15_X0/X13/M7_d N_X0/X13/13_X0/X13/M7_g
+ N_X0/X13/14_X0/X13/M7_s N_VDD_X0/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX0/X13/M8 N_VDD_X0/X13/M8_d N_B28_X0/X13/M8_g N_X0/X13/15_X0/X13/M8_s
+ N_VDD_X0/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X13/M9 N_X0/X13/15_X0/X13/M9_d N_A28_X0/X13/M9_g N_VDD_X0/X13/M9_s
+ N_VDD_X0/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X13/M10 N_VDD_X0/X13/M10_d N_X0/X13/14_X0/X13/M10_g N_X0/X13/16_X0/X13/M10_s
+ N_VDD_X0/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X13/M11 N_X0/X13/21_X0/X13/M11_d N_B28_X0/X13/M11_g N_VDD_X0/X13/M11_s
+ N_VDD_X0/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX0/X13/M12 N_X0/X13/13_X0/X13/M12_d N_A28_X0/X13/M12_g N_X0/X13/21_X0/X13/M12_s
+ N_VDD_X0/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X13/M13 N_VDD_X0/X13/M13_d N_X0/X13/13_X0/X13/M13_g N_X0/X13/17_X0/X13/M13_s
+ N_VDD_X0/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X13/X14/M0 N_GND_X0/X13/X14/M0_d N_X0/X13/18_X0/X13/X14/M0_g
+ N_SUM28_X0/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X13/X14/M1 N_X0/X13/X14/10_X0/X13/X14/M1_d N_X0/32_X0/X13/X14/M1_g
+ N_X0/X13/18_X0/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X13/X14/M2 N_GND_X0/X13/X14/M2_d N_3_X0/X13/X14/M2_g
+ N_X0/X13/X14/10_X0/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X13/X14/M3 N_X0/X13/X14/11_X0/X13/X14/M3_d N_X0/X13/16_X0/X13/X14/M3_g
+ N_GND_X0/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X13/X14/M4 N_X0/X13/18_X0/X13/X14/M4_d N_45_X0/X13/X14/M4_g
+ N_X0/X13/X14/11_X0/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X13/X14/M5 N_X0/X13/X14/9_X0/X13/X14/M5_d N_X0/X13/16_X0/X13/X14/M5_g
+ N_VDD_X0/X13/X14/M5_s N_VDD_X0/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X13/X14/M6 N_X0/X13/18_X0/X13/X14/M6_d N_X0/32_X0/X13/X14/M6_g
+ N_X0/X13/X14/9_X0/X13/X14/M6_s N_VDD_X0/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X14/M7 N_X0/X13/X14/9_X0/X13/X14/M7_d N_3_X0/X13/X14/M7_g
+ N_X0/X13/18_X0/X13/X14/M7_s N_VDD_X0/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X14/M8 N_VDD_X0/X13/X14/M8_d N_45_X0/X13/X14/M8_g
+ N_X0/X13/X14/9_X0/X13/X14/M8_s N_VDD_X0/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X13/X14/M9 N_VDD_X0/X13/X14/M9_d N_X0/X13/18_X0/X13/X14/M9_g
+ N_SUM28_X0/X13/X14/M9_s N_VDD_X0/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X13/X15/M0 N_GND_X0/X13/X15/M0_d N_X0/28_X0/X13/X15/M0_g
+ N_X0/37_X0/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X13/X15/M1 N_X0/X13/X15/10_X0/X13/X15/M1_d N_X0/X13/17_X0/X13/X15/M1_g
+ N_X0/28_X0/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX0/X13/X15/M2 N_GND_X0/X13/X15/M2_d N_45_X0/X13/X15/M2_g
+ N_X0/X13/X15/10_X0/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X13/X15/M3 N_X0/X13/X15/11_X0/X13/X15/M3_d N_B28_X0/X13/X15/M3_g
+ N_GND_X0/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X13/X15/M4 N_X0/28_X0/X13/X15/M4_d N_A28_X0/X13/X15/M4_g
+ N_X0/X13/X15/11_X0/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X13/X15/M5 N_X0/X13/X15/9_X0/X13/X15/M5_d N_B28_X0/X13/X15/M5_g
+ N_VDD_X0/X13/X15/M5_s N_VDD_X0/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X13/X15/M6 N_X0/28_X0/X13/X15/M6_d N_X0/X13/17_X0/X13/X15/M6_g
+ N_X0/X13/X15/9_X0/X13/X15/M6_s N_VDD_X0/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X15/M7 N_X0/X13/X15/9_X0/X13/X15/M7_d N_45_X0/X13/X15/M7_g
+ N_X0/28_X0/X13/X15/M7_s N_VDD_X0/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X15/M8 N_VDD_X0/X13/X15/M8_d N_A28_X0/X13/X15/M8_g
+ N_X0/X13/X15/9_X0/X13/X15/M8_s N_VDD_X0/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X13/X15/M9 N_VDD_X0/X13/X15/M9_d N_X0/28_X0/X13/X15/M9_g
+ N_X0/37_X0/X13/X15/M9_s N_VDD_X0/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X13/X16/M0 N_GND_X0/X13/X16/M0_d N_X0/X13/19_X0/X13/X16/M0_g
+ N_X0/32_X0/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X13/X16/M1 N_X0/X13/X16/10_X0/X13/X16/M1_d N_A28N_X0/X13/X16/M1_g
+ N_X0/X13/19_X0/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X13/X16/M2 N_GND_X0/X13/X16/M2_d N_B28_X0/X13/X16/M2_g
+ N_X0/X13/X16/10_X0/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X13/X16/M3 N_X0/X13/X16/11_X0/X13/X16/M3_d N_B28N_X0/X13/X16/M3_g
+ N_GND_X0/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X13/X16/M4 N_X0/X13/19_X0/X13/X16/M4_d N_A28_X0/X13/X16/M4_g
+ N_X0/X13/X16/11_X0/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X13/X16/M5 N_X0/X13/X16/9_X0/X13/X16/M5_d N_B28N_X0/X13/X16/M5_g
+ N_VDD_X0/X13/X16/M5_s N_VDD_X0/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X13/X16/M6 N_X0/X13/19_X0/X13/X16/M6_d N_A28N_X0/X13/X16/M6_g
+ N_X0/X13/X16/9_X0/X13/X16/M6_s N_VDD_X0/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X16/M7 N_X0/X13/X16/9_X0/X13/X16/M7_d N_B28_X0/X13/X16/M7_g
+ N_X0/X13/19_X0/X13/X16/M7_s N_VDD_X0/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X13/X16/M8 N_VDD_X0/X13/X16/M8_d N_A28_X0/X13/X16/M8_g
+ N_X0/X13/X16/9_X0/X13/X16/M8_s N_VDD_X0/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X13/X16/M9 N_VDD_X0/X13/X16/M9_d N_X0/X13/19_X0/X13/X16/M9_g
+ N_X0/32_X0/X13/X16/M9_s N_VDD_X0/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X14/M0 N_GND_X0/X14/M0_d N_X0/X14/14_X0/X14/M0_g N_X0/X14/16_X0/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X14/M1 N_GND_X0/X14/M1_d N_X0/X14/13_X0/X14/M1_g N_X0/X14/14_X0/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X14/M2 N_X0/X14/20_X0/X14/M2_d N_B31_X0/X14/M2_g N_GND_X0/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX0/X14/M3 N_X0/X14/14_X0/X14/M3_d N_A31_X0/X14/M3_g N_X0/X14/20_X0/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X14/M4 N_GND_X0/X14/M4_d N_X0/X14/13_X0/X14/M4_g N_X0/X14/17_X0/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X14/M5 N_X0/X14/13_X0/X14/M5_d N_B31_X0/X14/M5_g N_GND_X0/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX0/X14/M6 N_GND_X0/X14/M6_d N_A31_X0/X14/M6_g N_X0/X14/13_X0/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX0/X14/M7 N_X0/X14/15_X0/X14/M7_d N_X0/X14/13_X0/X14/M7_g
+ N_X0/X14/14_X0/X14/M7_s N_VDD_X0/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX0/X14/M8 N_VDD_X0/X14/M8_d N_B31_X0/X14/M8_g N_X0/X14/15_X0/X14/M8_s
+ N_VDD_X0/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX0/X14/M9 N_X0/X14/15_X0/X14/M9_d N_A31_X0/X14/M9_g N_VDD_X0/X14/M9_s
+ N_VDD_X0/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X14/M10 N_VDD_X0/X14/M10_d N_X0/X14/14_X0/X14/M10_g N_X0/X14/16_X0/X14/M10_s
+ N_VDD_X0/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X14/M11 N_X0/X14/21_X0/X14/M11_d N_B31_X0/X14/M11_g N_VDD_X0/X14/M11_s
+ N_VDD_X0/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX0/X14/M12 N_X0/X14/13_X0/X14/M12_d N_A31_X0/X14/M12_g N_X0/X14/21_X0/X14/M12_s
+ N_VDD_X0/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX0/X14/M13 N_VDD_X0/X14/M13_d N_X0/X14/13_X0/X14/M13_g N_X0/X14/17_X0/X14/M13_s
+ N_VDD_X0/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X14/X14/M0 N_GND_X0/X14/X14/M0_d N_X0/X14/18_X0/X14/X14/M0_g
+ N_SUM31_X0/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X14/X14/M1 N_X0/X14/X14/10_X0/X14/X14/M1_d N_X0/35_X0/X14/X14/M1_g
+ N_X0/X14/18_X0/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X14/X14/M2 N_GND_X0/X14/X14/M2_d N_X0/29_X0/X14/X14/M2_g
+ N_X0/X14/X14/10_X0/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X14/X14/M3 N_X0/X14/X14/11_X0/X14/X14/M3_d N_X0/X14/16_X0/X14/X14/M3_g
+ N_GND_X0/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X14/X14/M4 N_X0/X14/18_X0/X14/X14/M4_d N_X0/38_X0/X14/X14/M4_g
+ N_X0/X14/X14/11_X0/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X14/X14/M5 N_X0/X14/X14/9_X0/X14/X14/M5_d N_X0/X14/16_X0/X14/X14/M5_g
+ N_VDD_X0/X14/X14/M5_s N_VDD_X0/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X14/X14/M6 N_X0/X14/18_X0/X14/X14/M6_d N_X0/35_X0/X14/X14/M6_g
+ N_X0/X14/X14/9_X0/X14/X14/M6_s N_VDD_X0/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X14/M7 N_X0/X14/X14/9_X0/X14/X14/M7_d N_X0/29_X0/X14/X14/M7_g
+ N_X0/X14/18_X0/X14/X14/M7_s N_VDD_X0/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X14/M8 N_VDD_X0/X14/X14/M8_d N_X0/38_X0/X14/X14/M8_g
+ N_X0/X14/X14/9_X0/X14/X14/M8_s N_VDD_X0/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X14/X14/M9 N_VDD_X0/X14/X14/M9_d N_X0/X14/18_X0/X14/X14/M9_g
+ N_SUM31_X0/X14/X14/M9_s N_VDD_X0/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X14/X15/M0 N_GND_X0/X14/X15/M0_d N_X0/33_X0/X14/X15/M0_g
+ N_X0/34_X0/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X14/X15/M1 N_X0/X14/X15/10_X0/X14/X15/M1_d N_X0/X14/17_X0/X14/X15/M1_g
+ N_X0/33_X0/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX0/X14/X15/M2 N_GND_X0/X14/X15/M2_d N_X0/38_X0/X14/X15/M2_g
+ N_X0/X14/X15/10_X0/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X14/X15/M3 N_X0/X14/X15/11_X0/X14/X15/M3_d N_B31_X0/X14/X15/M3_g
+ N_GND_X0/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X14/X15/M4 N_X0/33_X0/X14/X15/M4_d N_A31_X0/X14/X15/M4_g
+ N_X0/X14/X15/11_X0/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X14/X15/M5 N_X0/X14/X15/9_X0/X14/X15/M5_d N_B31_X0/X14/X15/M5_g
+ N_VDD_X0/X14/X15/M5_s N_VDD_X0/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X14/X15/M6 N_X0/33_X0/X14/X15/M6_d N_X0/X14/17_X0/X14/X15/M6_g
+ N_X0/X14/X15/9_X0/X14/X15/M6_s N_VDD_X0/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X15/M7 N_X0/X14/X15/9_X0/X14/X15/M7_d N_X0/38_X0/X14/X15/M7_g
+ N_X0/33_X0/X14/X15/M7_s N_VDD_X0/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X15/M8 N_VDD_X0/X14/X15/M8_d N_A31_X0/X14/X15/M8_g
+ N_X0/X14/X15/9_X0/X14/X15/M8_s N_VDD_X0/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X14/X15/M9 N_VDD_X0/X14/X15/M9_d N_X0/33_X0/X14/X15/M9_g
+ N_X0/34_X0/X14/X15/M9_s N_VDD_X0/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX0/X14/X16/M0 N_GND_X0/X14/X16/M0_d N_X0/X14/19_X0/X14/X16/M0_g
+ N_X0/35_X0/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX0/X14/X16/M1 N_X0/X14/X16/10_X0/X14/X16/M1_d N_A31N_X0/X14/X16/M1_g
+ N_X0/X14/19_X0/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX0/X14/X16/M2 N_GND_X0/X14/X16/M2_d N_B31_X0/X14/X16/M2_g
+ N_X0/X14/X16/10_X0/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX0/X14/X16/M3 N_X0/X14/X16/11_X0/X14/X16/M3_d N_B31N_X0/X14/X16/M3_g
+ N_GND_X0/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX0/X14/X16/M4 N_X0/X14/19_X0/X14/X16/M4_d N_A31_X0/X14/X16/M4_g
+ N_X0/X14/X16/11_X0/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX0/X14/X16/M5 N_X0/X14/X16/9_X0/X14/X16/M5_d N_B31N_X0/X14/X16/M5_g
+ N_VDD_X0/X14/X16/M5_s N_VDD_X0/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX0/X14/X16/M6 N_X0/X14/19_X0/X14/X16/M6_d N_A31N_X0/X14/X16/M6_g
+ N_X0/X14/X16/9_X0/X14/X16/M6_s N_VDD_X0/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X16/M7 N_X0/X14/X16/9_X0/X14/X16/M7_d N_B31_X0/X14/X16/M7_g
+ N_X0/X14/19_X0/X14/X16/M7_s N_VDD_X0/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX0/X14/X16/M8 N_VDD_X0/X14/X16/M8_d N_A31_X0/X14/X16/M8_g
+ N_X0/X14/X16/9_X0/X14/X16/M8_s N_VDD_X0/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX0/X14/X16/M9 N_VDD_X0/X14/X16/M9_d N_X0/X14/19_X0/X14/X16/M9_g
+ N_X0/35_X0/X14/X16/M9_s N_VDD_X0/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/M0 N_GND_X1/M0_d N_X1/39_X1/M0_g N_X1/40_X1/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/M1 N_X1/41_X1/M1_d N_X1/32_X1/M1_g N_GND_X1/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX1/M2 N_X1/42_X1/M2_d N_X1/31_X1/M2_g N_X1/41_X1/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX1/M3 N_X1/43_X1/M3_d N_X1/30_X1/M3_g N_X1/42_X1/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX1/M4 N_X1/39_X1/M4_d N_X1/35_X1/M4_g N_X1/43_X1/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX1/M5 N_VDD_X1/M5_d N_X1/39_X1/M5_g N_X1/40_X1/M5_s N_VDD_X1/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/M6 N_X1/39_X1/M6_d N_X1/32_X1/M6_g N_VDD_X1/M6_s N_VDD_X1/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX1/M7 N_VDD_X1/M7_d N_X1/31_X1/M7_g N_X1/39_X1/M7_s N_VDD_X1/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX1/M8 N_X1/39_X1/M8_d N_X1/30_X1/M8_g N_VDD_X1/M8_s N_VDD_X1/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX1/M9 N_VDD_X1/M9_d N_X1/35_X1/M9_g N_X1/39_X1/M9_s N_VDD_X1/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX1/X10/M0 N_GND_X1/X10/M0_d N_3_X1/X10/M0_g N_45_X1/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X10/M1 N_X1/X10/10_X1/X10/M1_d N_46_X1/X10/M1_g N_3_X1/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X10/M2 N_GND_X1/X10/M2_d N_X1/40_X1/X10/M2_g N_X1/X10/10_X1/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X10/M3 N_X1/X10/11_X1/X10/M3_d N_X1/39_X1/X10/M3_g N_GND_X1/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X10/M4 N_3_X1/X10/M4_d N_X1/34_X1/X10/M4_g N_X1/X10/11_X1/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X10/M5 N_X1/X10/9_X1/X10/M5_d N_X1/39_X1/X10/M5_g N_VDD_X1/X10/M5_s
+ N_VDD_X1/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX1/X10/M6 N_3_X1/X10/M6_d N_46_X1/X10/M6_g N_X1/X10/9_X1/X10/M6_s
+ N_VDD_X1/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X10/M7 N_X1/X10/9_X1/X10/M7_d N_X1/40_X1/X10/M7_g N_3_X1/X10/M7_s
+ N_VDD_X1/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X10/M8 N_VDD_X1/X10/M8_d N_X1/34_X1/X10/M8_g N_X1/X10/9_X1/X10/M8_s
+ N_VDD_X1/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X10/M9 N_VDD_X1/X10/M9_d N_3_X1/X10/M9_g N_45_X1/X10/M9_s N_VDD_X1/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X11/M0 N_GND_X1/X11/M0_d N_X1/X11/14_X1/X11/M0_g N_X1/X11/16_X1/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X11/M1 N_GND_X1/X11/M1_d N_X1/X11/13_X1/X11/M1_g N_X1/X11/14_X1/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X11/M2 N_X1/X11/20_X1/X11/M2_d N_B26_X1/X11/M2_g N_GND_X1/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X11/M3 N_X1/X11/14_X1/X11/M3_d N_A26_X1/X11/M3_g N_X1/X11/20_X1/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X11/M4 N_GND_X1/X11/M4_d N_X1/X11/13_X1/X11/M4_g N_X1/X11/17_X1/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X11/M5 N_X1/X11/13_X1/X11/M5_d N_B26_X1/X11/M5_g N_GND_X1/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X11/M6 N_GND_X1/X11/M6_d N_A26_X1/X11/M6_g N_X1/X11/13_X1/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X11/M7 N_X1/X11/15_X1/X11/M7_d N_X1/X11/13_X1/X11/M7_g
+ N_X1/X11/14_X1/X11/M7_s N_VDD_X1/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX1/X11/M8 N_VDD_X1/X11/M8_d N_B26_X1/X11/M8_g N_X1/X11/15_X1/X11/M8_s
+ N_VDD_X1/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X11/M9 N_X1/X11/15_X1/X11/M9_d N_A26_X1/X11/M9_g N_VDD_X1/X11/M9_s
+ N_VDD_X1/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X11/M10 N_VDD_X1/X11/M10_d N_X1/X11/14_X1/X11/M10_g N_X1/X11/16_X1/X11/M10_s
+ N_VDD_X1/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X11/M11 N_X1/X11/21_X1/X11/M11_d N_B26_X1/X11/M11_g N_VDD_X1/X11/M11_s
+ N_VDD_X1/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX1/X11/M12 N_X1/X11/13_X1/X11/M12_d N_A26_X1/X11/M12_g N_X1/X11/21_X1/X11/M12_s
+ N_VDD_X1/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X11/M13 N_VDD_X1/X11/M13_d N_X1/X11/13_X1/X11/M13_g N_X1/X11/17_X1/X11/M13_s
+ N_VDD_X1/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X11/X14/M0 N_GND_X1/X11/X14/M0_d N_X1/X11/18_X1/X11/X14/M0_g
+ N_SUM26_X1/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X11/X14/M1 N_X1/X11/X14/10_X1/X11/X14/M1_d N_X1/30_X1/X11/X14/M1_g
+ N_X1/X11/18_X1/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X11/X14/M2 N_GND_X1/X11/X14/M2_d N_X1/27_X1/X11/X14/M2_g
+ N_X1/X11/X14/10_X1/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X11/X14/M3 N_X1/X11/X14/11_X1/X11/X14/M3_d N_X1/X11/16_X1/X11/X14/M3_g
+ N_GND_X1/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X11/X14/M4 N_X1/X11/18_X1/X11/X14/M4_d N_X1/36_X1/X11/X14/M4_g
+ N_X1/X11/X14/11_X1/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X11/X14/M5 N_X1/X11/X14/9_X1/X11/X14/M5_d N_X1/X11/16_X1/X11/X14/M5_g
+ N_VDD_X1/X11/X14/M5_s N_VDD_X1/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X11/X14/M6 N_X1/X11/18_X1/X11/X14/M6_d N_X1/30_X1/X11/X14/M6_g
+ N_X1/X11/X14/9_X1/X11/X14/M6_s N_VDD_X1/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X14/M7 N_X1/X11/X14/9_X1/X11/X14/M7_d N_X1/27_X1/X11/X14/M7_g
+ N_X1/X11/18_X1/X11/X14/M7_s N_VDD_X1/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X14/M8 N_VDD_X1/X11/X14/M8_d N_X1/36_X1/X11/X14/M8_g
+ N_X1/X11/X14/9_X1/X11/X14/M8_s N_VDD_X1/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X11/X14/M9 N_VDD_X1/X11/X14/M9_d N_X1/X11/18_X1/X11/X14/M9_g
+ N_SUM26_X1/X11/X14/M9_s N_VDD_X1/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X11/X15/M0 N_GND_X1/X11/X15/M0_d N_X1/29_X1/X11/X15/M0_g
+ N_X1/38_X1/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X11/X15/M1 N_X1/X11/X15/10_X1/X11/X15/M1_d N_X1/X11/17_X1/X11/X15/M1_g
+ N_X1/29_X1/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX1/X11/X15/M2 N_GND_X1/X11/X15/M2_d N_X1/36_X1/X11/X15/M2_g
+ N_X1/X11/X15/10_X1/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X11/X15/M3 N_X1/X11/X15/11_X1/X11/X15/M3_d N_B26_X1/X11/X15/M3_g
+ N_GND_X1/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X11/X15/M4 N_X1/29_X1/X11/X15/M4_d N_A26_X1/X11/X15/M4_g
+ N_X1/X11/X15/11_X1/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X11/X15/M5 N_X1/X11/X15/9_X1/X11/X15/M5_d N_B26_X1/X11/X15/M5_g
+ N_VDD_X1/X11/X15/M5_s N_VDD_X1/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X11/X15/M6 N_X1/29_X1/X11/X15/M6_d N_X1/X11/17_X1/X11/X15/M6_g
+ N_X1/X11/X15/9_X1/X11/X15/M6_s N_VDD_X1/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X15/M7 N_X1/X11/X15/9_X1/X11/X15/M7_d N_X1/36_X1/X11/X15/M7_g
+ N_X1/29_X1/X11/X15/M7_s N_VDD_X1/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X15/M8 N_VDD_X1/X11/X15/M8_d N_A26_X1/X11/X15/M8_g
+ N_X1/X11/X15/9_X1/X11/X15/M8_s N_VDD_X1/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X11/X15/M9 N_VDD_X1/X11/X15/M9_d N_X1/29_X1/X11/X15/M9_g
+ N_X1/38_X1/X11/X15/M9_s N_VDD_X1/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X11/X16/M0 N_GND_X1/X11/X16/M0_d N_X1/X11/19_X1/X11/X16/M0_g
+ N_X1/30_X1/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X11/X16/M1 N_X1/X11/X16/10_X1/X11/X16/M1_d N_A26N_X1/X11/X16/M1_g
+ N_X1/X11/19_X1/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X11/X16/M2 N_GND_X1/X11/X16/M2_d N_B26_X1/X11/X16/M2_g
+ N_X1/X11/X16/10_X1/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X11/X16/M3 N_X1/X11/X16/11_X1/X11/X16/M3_d N_B26N_X1/X11/X16/M3_g
+ N_GND_X1/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X11/X16/M4 N_X1/X11/19_X1/X11/X16/M4_d N_A26_X1/X11/X16/M4_g
+ N_X1/X11/X16/11_X1/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X11/X16/M5 N_X1/X11/X16/9_X1/X11/X16/M5_d N_B26N_X1/X11/X16/M5_g
+ N_VDD_X1/X11/X16/M5_s N_VDD_X1/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X11/X16/M6 N_X1/X11/19_X1/X11/X16/M6_d N_A26N_X1/X11/X16/M6_g
+ N_X1/X11/X16/9_X1/X11/X16/M6_s N_VDD_X1/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X16/M7 N_X1/X11/X16/9_X1/X11/X16/M7_d N_B26_X1/X11/X16/M7_g
+ N_X1/X11/19_X1/X11/X16/M7_s N_VDD_X1/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X11/X16/M8 N_VDD_X1/X11/X16/M8_d N_A26_X1/X11/X16/M8_g
+ N_X1/X11/X16/9_X1/X11/X16/M8_s N_VDD_X1/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X11/X16/M9 N_VDD_X1/X11/X16/M9_d N_X1/X11/19_X1/X11/X16/M9_g
+ N_X1/30_X1/X11/X16/M9_s N_VDD_X1/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X12/M0 N_GND_X1/X12/M0_d N_X1/X12/14_X1/X12/M0_g N_X1/X12/16_X1/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X12/M1 N_GND_X1/X12/M1_d N_X1/X12/13_X1/X12/M1_g N_X1/X12/14_X1/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X12/M2 N_X1/X12/20_X1/X12/M2_d N_B25_X1/X12/M2_g N_GND_X1/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X12/M3 N_X1/X12/14_X1/X12/M3_d N_A25_X1/X12/M3_g N_X1/X12/20_X1/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X12/M4 N_GND_X1/X12/M4_d N_X1/X12/13_X1/X12/M4_g N_X1/X12/17_X1/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X12/M5 N_X1/X12/13_X1/X12/M5_d N_B25_X1/X12/M5_g N_GND_X1/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X12/M6 N_GND_X1/X12/M6_d N_A25_X1/X12/M6_g N_X1/X12/13_X1/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X12/M7 N_X1/X12/15_X1/X12/M7_d N_X1/X12/13_X1/X12/M7_g
+ N_X1/X12/14_X1/X12/M7_s N_VDD_X1/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX1/X12/M8 N_VDD_X1/X12/M8_d N_B25_X1/X12/M8_g N_X1/X12/15_X1/X12/M8_s
+ N_VDD_X1/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X12/M9 N_X1/X12/15_X1/X12/M9_d N_A25_X1/X12/M9_g N_VDD_X1/X12/M9_s
+ N_VDD_X1/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X12/M10 N_VDD_X1/X12/M10_d N_X1/X12/14_X1/X12/M10_g N_X1/X12/16_X1/X12/M10_s
+ N_VDD_X1/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X12/M11 N_X1/X12/21_X1/X12/M11_d N_B25_X1/X12/M11_g N_VDD_X1/X12/M11_s
+ N_VDD_X1/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX1/X12/M12 N_X1/X12/13_X1/X12/M12_d N_A25_X1/X12/M12_g N_X1/X12/21_X1/X12/M12_s
+ N_VDD_X1/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X12/M13 N_VDD_X1/X12/M13_d N_X1/X12/13_X1/X12/M13_g N_X1/X12/17_X1/X12/M13_s
+ N_VDD_X1/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X12/X14/M0 N_GND_X1/X12/X14/M0_d N_X1/X12/18_X1/X12/X14/M0_g
+ N_SUM25_X1/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X12/X14/M1 N_X1/X12/X14/10_X1/X12/X14/M1_d N_X1/31_X1/X12/X14/M1_g
+ N_X1/X12/18_X1/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X12/X14/M2 N_GND_X1/X12/X14/M2_d N_X1/28_X1/X12/X14/M2_g
+ N_X1/X12/X14/10_X1/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X12/X14/M3 N_X1/X12/X14/11_X1/X12/X14/M3_d N_X1/X12/16_X1/X12/X14/M3_g
+ N_GND_X1/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X12/X14/M4 N_X1/X12/18_X1/X12/X14/M4_d N_X1/37_X1/X12/X14/M4_g
+ N_X1/X12/X14/11_X1/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X12/X14/M5 N_X1/X12/X14/9_X1/X12/X14/M5_d N_X1/X12/16_X1/X12/X14/M5_g
+ N_VDD_X1/X12/X14/M5_s N_VDD_X1/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X12/X14/M6 N_X1/X12/18_X1/X12/X14/M6_d N_X1/31_X1/X12/X14/M6_g
+ N_X1/X12/X14/9_X1/X12/X14/M6_s N_VDD_X1/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X14/M7 N_X1/X12/X14/9_X1/X12/X14/M7_d N_X1/28_X1/X12/X14/M7_g
+ N_X1/X12/18_X1/X12/X14/M7_s N_VDD_X1/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X14/M8 N_VDD_X1/X12/X14/M8_d N_X1/37_X1/X12/X14/M8_g
+ N_X1/X12/X14/9_X1/X12/X14/M8_s N_VDD_X1/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X12/X14/M9 N_VDD_X1/X12/X14/M9_d N_X1/X12/18_X1/X12/X14/M9_g
+ N_SUM25_X1/X12/X14/M9_s N_VDD_X1/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X12/X15/M0 N_GND_X1/X12/X15/M0_d N_X1/27_X1/X12/X15/M0_g
+ N_X1/36_X1/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X12/X15/M1 N_X1/X12/X15/10_X1/X12/X15/M1_d N_X1/X12/17_X1/X12/X15/M1_g
+ N_X1/27_X1/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX1/X12/X15/M2 N_GND_X1/X12/X15/M2_d N_X1/37_X1/X12/X15/M2_g
+ N_X1/X12/X15/10_X1/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X12/X15/M3 N_X1/X12/X15/11_X1/X12/X15/M3_d N_B25_X1/X12/X15/M3_g
+ N_GND_X1/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X12/X15/M4 N_X1/27_X1/X12/X15/M4_d N_A25_X1/X12/X15/M4_g
+ N_X1/X12/X15/11_X1/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X12/X15/M5 N_X1/X12/X15/9_X1/X12/X15/M5_d N_B25_X1/X12/X15/M5_g
+ N_VDD_X1/X12/X15/M5_s N_VDD_X1/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X12/X15/M6 N_X1/27_X1/X12/X15/M6_d N_X1/X12/17_X1/X12/X15/M6_g
+ N_X1/X12/X15/9_X1/X12/X15/M6_s N_VDD_X1/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X15/M7 N_X1/X12/X15/9_X1/X12/X15/M7_d N_X1/37_X1/X12/X15/M7_g
+ N_X1/27_X1/X12/X15/M7_s N_VDD_X1/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X15/M8 N_VDD_X1/X12/X15/M8_d N_A25_X1/X12/X15/M8_g
+ N_X1/X12/X15/9_X1/X12/X15/M8_s N_VDD_X1/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X12/X15/M9 N_VDD_X1/X12/X15/M9_d N_X1/27_X1/X12/X15/M9_g
+ N_X1/36_X1/X12/X15/M9_s N_VDD_X1/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X12/X16/M0 N_GND_X1/X12/X16/M0_d N_X1/X12/19_X1/X12/X16/M0_g
+ N_X1/31_X1/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X12/X16/M1 N_X1/X12/X16/10_X1/X12/X16/M1_d N_A25N_X1/X12/X16/M1_g
+ N_X1/X12/19_X1/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X12/X16/M2 N_GND_X1/X12/X16/M2_d N_B25_X1/X12/X16/M2_g
+ N_X1/X12/X16/10_X1/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X12/X16/M3 N_X1/X12/X16/11_X1/X12/X16/M3_d N_B25N_X1/X12/X16/M3_g
+ N_GND_X1/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X12/X16/M4 N_X1/X12/19_X1/X12/X16/M4_d N_A25_X1/X12/X16/M4_g
+ N_X1/X12/X16/11_X1/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X12/X16/M5 N_X1/X12/X16/9_X1/X12/X16/M5_d N_B25N_X1/X12/X16/M5_g
+ N_VDD_X1/X12/X16/M5_s N_VDD_X1/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X12/X16/M6 N_X1/X12/19_X1/X12/X16/M6_d N_A25N_X1/X12/X16/M6_g
+ N_X1/X12/X16/9_X1/X12/X16/M6_s N_VDD_X1/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X16/M7 N_X1/X12/X16/9_X1/X12/X16/M7_d N_B25_X1/X12/X16/M7_g
+ N_X1/X12/19_X1/X12/X16/M7_s N_VDD_X1/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X12/X16/M8 N_VDD_X1/X12/X16/M8_d N_A25_X1/X12/X16/M8_g
+ N_X1/X12/X16/9_X1/X12/X16/M8_s N_VDD_X1/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X12/X16/M9 N_VDD_X1/X12/X16/M9_d N_X1/X12/19_X1/X12/X16/M9_g
+ N_X1/31_X1/X12/X16/M9_s N_VDD_X1/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X13/M0 N_GND_X1/X13/M0_d N_X1/X13/14_X1/X13/M0_g N_X1/X13/16_X1/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X13/M1 N_GND_X1/X13/M1_d N_X1/X13/13_X1/X13/M1_g N_X1/X13/14_X1/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X13/M2 N_X1/X13/20_X1/X13/M2_d N_B24_X1/X13/M2_g N_GND_X1/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X13/M3 N_X1/X13/14_X1/X13/M3_d N_A24_X1/X13/M3_g N_X1/X13/20_X1/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X13/M4 N_GND_X1/X13/M4_d N_X1/X13/13_X1/X13/M4_g N_X1/X13/17_X1/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X13/M5 N_X1/X13/13_X1/X13/M5_d N_B24_X1/X13/M5_g N_GND_X1/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X13/M6 N_GND_X1/X13/M6_d N_A24_X1/X13/M6_g N_X1/X13/13_X1/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X13/M7 N_X1/X13/15_X1/X13/M7_d N_X1/X13/13_X1/X13/M7_g
+ N_X1/X13/14_X1/X13/M7_s N_VDD_X1/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX1/X13/M8 N_VDD_X1/X13/M8_d N_B24_X1/X13/M8_g N_X1/X13/15_X1/X13/M8_s
+ N_VDD_X1/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X13/M9 N_X1/X13/15_X1/X13/M9_d N_A24_X1/X13/M9_g N_VDD_X1/X13/M9_s
+ N_VDD_X1/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X13/M10 N_VDD_X1/X13/M10_d N_X1/X13/14_X1/X13/M10_g N_X1/X13/16_X1/X13/M10_s
+ N_VDD_X1/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X13/M11 N_X1/X13/21_X1/X13/M11_d N_B24_X1/X13/M11_g N_VDD_X1/X13/M11_s
+ N_VDD_X1/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX1/X13/M12 N_X1/X13/13_X1/X13/M12_d N_A24_X1/X13/M12_g N_X1/X13/21_X1/X13/M12_s
+ N_VDD_X1/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X13/M13 N_VDD_X1/X13/M13_d N_X1/X13/13_X1/X13/M13_g N_X1/X13/17_X1/X13/M13_s
+ N_VDD_X1/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X13/X14/M0 N_GND_X1/X13/X14/M0_d N_X1/X13/18_X1/X13/X14/M0_g
+ N_SUM24_X1/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X13/X14/M1 N_X1/X13/X14/10_X1/X13/X14/M1_d N_X1/32_X1/X13/X14/M1_g
+ N_X1/X13/18_X1/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X13/X14/M2 N_GND_X1/X13/X14/M2_d N_4_X1/X13/X14/M2_g
+ N_X1/X13/X14/10_X1/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X13/X14/M3 N_X1/X13/X14/11_X1/X13/X14/M3_d N_X1/X13/16_X1/X13/X14/M3_g
+ N_GND_X1/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X13/X14/M4 N_X1/X13/18_X1/X13/X14/M4_d N_46_X1/X13/X14/M4_g
+ N_X1/X13/X14/11_X1/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X13/X14/M5 N_X1/X13/X14/9_X1/X13/X14/M5_d N_X1/X13/16_X1/X13/X14/M5_g
+ N_VDD_X1/X13/X14/M5_s N_VDD_X1/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X13/X14/M6 N_X1/X13/18_X1/X13/X14/M6_d N_X1/32_X1/X13/X14/M6_g
+ N_X1/X13/X14/9_X1/X13/X14/M6_s N_VDD_X1/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X14/M7 N_X1/X13/X14/9_X1/X13/X14/M7_d N_4_X1/X13/X14/M7_g
+ N_X1/X13/18_X1/X13/X14/M7_s N_VDD_X1/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X14/M8 N_VDD_X1/X13/X14/M8_d N_46_X1/X13/X14/M8_g
+ N_X1/X13/X14/9_X1/X13/X14/M8_s N_VDD_X1/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X13/X14/M9 N_VDD_X1/X13/X14/M9_d N_X1/X13/18_X1/X13/X14/M9_g
+ N_SUM24_X1/X13/X14/M9_s N_VDD_X1/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X13/X15/M0 N_GND_X1/X13/X15/M0_d N_X1/28_X1/X13/X15/M0_g
+ N_X1/37_X1/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X13/X15/M1 N_X1/X13/X15/10_X1/X13/X15/M1_d N_X1/X13/17_X1/X13/X15/M1_g
+ N_X1/28_X1/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX1/X13/X15/M2 N_GND_X1/X13/X15/M2_d N_46_X1/X13/X15/M2_g
+ N_X1/X13/X15/10_X1/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X13/X15/M3 N_X1/X13/X15/11_X1/X13/X15/M3_d N_B24_X1/X13/X15/M3_g
+ N_GND_X1/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X13/X15/M4 N_X1/28_X1/X13/X15/M4_d N_A24_X1/X13/X15/M4_g
+ N_X1/X13/X15/11_X1/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X13/X15/M5 N_X1/X13/X15/9_X1/X13/X15/M5_d N_B24_X1/X13/X15/M5_g
+ N_VDD_X1/X13/X15/M5_s N_VDD_X1/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X13/X15/M6 N_X1/28_X1/X13/X15/M6_d N_X1/X13/17_X1/X13/X15/M6_g
+ N_X1/X13/X15/9_X1/X13/X15/M6_s N_VDD_X1/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X15/M7 N_X1/X13/X15/9_X1/X13/X15/M7_d N_46_X1/X13/X15/M7_g
+ N_X1/28_X1/X13/X15/M7_s N_VDD_X1/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X15/M8 N_VDD_X1/X13/X15/M8_d N_A24_X1/X13/X15/M8_g
+ N_X1/X13/X15/9_X1/X13/X15/M8_s N_VDD_X1/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X13/X15/M9 N_VDD_X1/X13/X15/M9_d N_X1/28_X1/X13/X15/M9_g
+ N_X1/37_X1/X13/X15/M9_s N_VDD_X1/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X13/X16/M0 N_GND_X1/X13/X16/M0_d N_X1/X13/19_X1/X13/X16/M0_g
+ N_X1/32_X1/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X13/X16/M1 N_X1/X13/X16/10_X1/X13/X16/M1_d N_A24N_X1/X13/X16/M1_g
+ N_X1/X13/19_X1/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X13/X16/M2 N_GND_X1/X13/X16/M2_d N_B24_X1/X13/X16/M2_g
+ N_X1/X13/X16/10_X1/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X13/X16/M3 N_X1/X13/X16/11_X1/X13/X16/M3_d N_B24N_X1/X13/X16/M3_g
+ N_GND_X1/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X13/X16/M4 N_X1/X13/19_X1/X13/X16/M4_d N_A24_X1/X13/X16/M4_g
+ N_X1/X13/X16/11_X1/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X13/X16/M5 N_X1/X13/X16/9_X1/X13/X16/M5_d N_B24N_X1/X13/X16/M5_g
+ N_VDD_X1/X13/X16/M5_s N_VDD_X1/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X13/X16/M6 N_X1/X13/19_X1/X13/X16/M6_d N_A24N_X1/X13/X16/M6_g
+ N_X1/X13/X16/9_X1/X13/X16/M6_s N_VDD_X1/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X16/M7 N_X1/X13/X16/9_X1/X13/X16/M7_d N_B24_X1/X13/X16/M7_g
+ N_X1/X13/19_X1/X13/X16/M7_s N_VDD_X1/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X13/X16/M8 N_VDD_X1/X13/X16/M8_d N_A24_X1/X13/X16/M8_g
+ N_X1/X13/X16/9_X1/X13/X16/M8_s N_VDD_X1/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X13/X16/M9 N_VDD_X1/X13/X16/M9_d N_X1/X13/19_X1/X13/X16/M9_g
+ N_X1/32_X1/X13/X16/M9_s N_VDD_X1/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X14/M0 N_GND_X1/X14/M0_d N_X1/X14/14_X1/X14/M0_g N_X1/X14/16_X1/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X14/M1 N_GND_X1/X14/M1_d N_X1/X14/13_X1/X14/M1_g N_X1/X14/14_X1/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X14/M2 N_X1/X14/20_X1/X14/M2_d N_B27_X1/X14/M2_g N_GND_X1/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX1/X14/M3 N_X1/X14/14_X1/X14/M3_d N_A27_X1/X14/M3_g N_X1/X14/20_X1/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X14/M4 N_GND_X1/X14/M4_d N_X1/X14/13_X1/X14/M4_g N_X1/X14/17_X1/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X14/M5 N_X1/X14/13_X1/X14/M5_d N_B27_X1/X14/M5_g N_GND_X1/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX1/X14/M6 N_GND_X1/X14/M6_d N_A27_X1/X14/M6_g N_X1/X14/13_X1/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX1/X14/M7 N_X1/X14/15_X1/X14/M7_d N_X1/X14/13_X1/X14/M7_g
+ N_X1/X14/14_X1/X14/M7_s N_VDD_X1/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX1/X14/M8 N_VDD_X1/X14/M8_d N_B27_X1/X14/M8_g N_X1/X14/15_X1/X14/M8_s
+ N_VDD_X1/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX1/X14/M9 N_X1/X14/15_X1/X14/M9_d N_A27_X1/X14/M9_g N_VDD_X1/X14/M9_s
+ N_VDD_X1/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X14/M10 N_VDD_X1/X14/M10_d N_X1/X14/14_X1/X14/M10_g N_X1/X14/16_X1/X14/M10_s
+ N_VDD_X1/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X14/M11 N_X1/X14/21_X1/X14/M11_d N_B27_X1/X14/M11_g N_VDD_X1/X14/M11_s
+ N_VDD_X1/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX1/X14/M12 N_X1/X14/13_X1/X14/M12_d N_A27_X1/X14/M12_g N_X1/X14/21_X1/X14/M12_s
+ N_VDD_X1/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX1/X14/M13 N_VDD_X1/X14/M13_d N_X1/X14/13_X1/X14/M13_g N_X1/X14/17_X1/X14/M13_s
+ N_VDD_X1/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X14/X14/M0 N_GND_X1/X14/X14/M0_d N_X1/X14/18_X1/X14/X14/M0_g
+ N_SUM27_X1/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X14/X14/M1 N_X1/X14/X14/10_X1/X14/X14/M1_d N_X1/35_X1/X14/X14/M1_g
+ N_X1/X14/18_X1/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X14/X14/M2 N_GND_X1/X14/X14/M2_d N_X1/29_X1/X14/X14/M2_g
+ N_X1/X14/X14/10_X1/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X14/X14/M3 N_X1/X14/X14/11_X1/X14/X14/M3_d N_X1/X14/16_X1/X14/X14/M3_g
+ N_GND_X1/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X14/X14/M4 N_X1/X14/18_X1/X14/X14/M4_d N_X1/38_X1/X14/X14/M4_g
+ N_X1/X14/X14/11_X1/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X14/X14/M5 N_X1/X14/X14/9_X1/X14/X14/M5_d N_X1/X14/16_X1/X14/X14/M5_g
+ N_VDD_X1/X14/X14/M5_s N_VDD_X1/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X14/X14/M6 N_X1/X14/18_X1/X14/X14/M6_d N_X1/35_X1/X14/X14/M6_g
+ N_X1/X14/X14/9_X1/X14/X14/M6_s N_VDD_X1/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X14/M7 N_X1/X14/X14/9_X1/X14/X14/M7_d N_X1/29_X1/X14/X14/M7_g
+ N_X1/X14/18_X1/X14/X14/M7_s N_VDD_X1/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X14/M8 N_VDD_X1/X14/X14/M8_d N_X1/38_X1/X14/X14/M8_g
+ N_X1/X14/X14/9_X1/X14/X14/M8_s N_VDD_X1/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X14/X14/M9 N_VDD_X1/X14/X14/M9_d N_X1/X14/18_X1/X14/X14/M9_g
+ N_SUM27_X1/X14/X14/M9_s N_VDD_X1/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X14/X15/M0 N_GND_X1/X14/X15/M0_d N_X1/33_X1/X14/X15/M0_g
+ N_X1/34_X1/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X14/X15/M1 N_X1/X14/X15/10_X1/X14/X15/M1_d N_X1/X14/17_X1/X14/X15/M1_g
+ N_X1/33_X1/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX1/X14/X15/M2 N_GND_X1/X14/X15/M2_d N_X1/38_X1/X14/X15/M2_g
+ N_X1/X14/X15/10_X1/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X14/X15/M3 N_X1/X14/X15/11_X1/X14/X15/M3_d N_B27_X1/X14/X15/M3_g
+ N_GND_X1/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X14/X15/M4 N_X1/33_X1/X14/X15/M4_d N_A27_X1/X14/X15/M4_g
+ N_X1/X14/X15/11_X1/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X14/X15/M5 N_X1/X14/X15/9_X1/X14/X15/M5_d N_B27_X1/X14/X15/M5_g
+ N_VDD_X1/X14/X15/M5_s N_VDD_X1/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X14/X15/M6 N_X1/33_X1/X14/X15/M6_d N_X1/X14/17_X1/X14/X15/M6_g
+ N_X1/X14/X15/9_X1/X14/X15/M6_s N_VDD_X1/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X15/M7 N_X1/X14/X15/9_X1/X14/X15/M7_d N_X1/38_X1/X14/X15/M7_g
+ N_X1/33_X1/X14/X15/M7_s N_VDD_X1/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X15/M8 N_VDD_X1/X14/X15/M8_d N_A27_X1/X14/X15/M8_g
+ N_X1/X14/X15/9_X1/X14/X15/M8_s N_VDD_X1/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X14/X15/M9 N_VDD_X1/X14/X15/M9_d N_X1/33_X1/X14/X15/M9_g
+ N_X1/34_X1/X14/X15/M9_s N_VDD_X1/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX1/X14/X16/M0 N_GND_X1/X14/X16/M0_d N_X1/X14/19_X1/X14/X16/M0_g
+ N_X1/35_X1/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX1/X14/X16/M1 N_X1/X14/X16/10_X1/X14/X16/M1_d N_A27N_X1/X14/X16/M1_g
+ N_X1/X14/19_X1/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX1/X14/X16/M2 N_GND_X1/X14/X16/M2_d N_B27_X1/X14/X16/M2_g
+ N_X1/X14/X16/10_X1/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX1/X14/X16/M3 N_X1/X14/X16/11_X1/X14/X16/M3_d N_B27N_X1/X14/X16/M3_g
+ N_GND_X1/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX1/X14/X16/M4 N_X1/X14/19_X1/X14/X16/M4_d N_A27_X1/X14/X16/M4_g
+ N_X1/X14/X16/11_X1/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX1/X14/X16/M5 N_X1/X14/X16/9_X1/X14/X16/M5_d N_B27N_X1/X14/X16/M5_g
+ N_VDD_X1/X14/X16/M5_s N_VDD_X1/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX1/X14/X16/M6 N_X1/X14/19_X1/X14/X16/M6_d N_A27N_X1/X14/X16/M6_g
+ N_X1/X14/X16/9_X1/X14/X16/M6_s N_VDD_X1/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X16/M7 N_X1/X14/X16/9_X1/X14/X16/M7_d N_B27_X1/X14/X16/M7_g
+ N_X1/X14/19_X1/X14/X16/M7_s N_VDD_X1/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX1/X14/X16/M8 N_VDD_X1/X14/X16/M8_d N_A27_X1/X14/X16/M8_g
+ N_X1/X14/X16/9_X1/X14/X16/M8_s N_VDD_X1/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX1/X14/X16/M9 N_VDD_X1/X14/X16/M9_d N_X1/X14/19_X1/X14/X16/M9_g
+ N_X1/35_X1/X14/X16/M9_s N_VDD_X1/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/M0 N_GND_X2/M0_d N_X2/39_X2/M0_g N_X2/40_X2/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/M1 N_X2/41_X2/M1_d N_X2/32_X2/M1_g N_GND_X2/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX2/M2 N_X2/42_X2/M2_d N_X2/31_X2/M2_g N_X2/41_X2/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX2/M3 N_X2/43_X2/M3_d N_X2/30_X2/M3_g N_X2/42_X2/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX2/M4 N_X2/39_X2/M4_d N_X2/35_X2/M4_g N_X2/43_X2/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX2/M5 N_VDD_X2/M5_d N_X2/39_X2/M5_g N_X2/40_X2/M5_s N_VDD_X2/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/M6 N_X2/39_X2/M6_d N_X2/32_X2/M6_g N_VDD_X2/M6_s N_VDD_X2/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX2/M7 N_VDD_X2/M7_d N_X2/31_X2/M7_g N_X2/39_X2/M7_s N_VDD_X2/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX2/M8 N_X2/39_X2/M8_d N_X2/30_X2/M8_g N_VDD_X2/M8_s N_VDD_X2/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX2/M9 N_VDD_X2/M9_d N_X2/35_X2/M9_g N_X2/39_X2/M9_s N_VDD_X2/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX2/X10/M0 N_GND_X2/X10/M0_d N_4_X2/X10/M0_g N_46_X2/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X10/M1 N_X2/X10/10_X2/X10/M1_d N_47_X2/X10/M1_g N_4_X2/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X10/M2 N_GND_X2/X10/M2_d N_X2/40_X2/X10/M2_g N_X2/X10/10_X2/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X10/M3 N_X2/X10/11_X2/X10/M3_d N_X2/39_X2/X10/M3_g N_GND_X2/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X10/M4 N_4_X2/X10/M4_d N_X2/34_X2/X10/M4_g N_X2/X10/11_X2/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X10/M5 N_X2/X10/9_X2/X10/M5_d N_X2/39_X2/X10/M5_g N_VDD_X2/X10/M5_s
+ N_VDD_X2/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX2/X10/M6 N_4_X2/X10/M6_d N_47_X2/X10/M6_g N_X2/X10/9_X2/X10/M6_s
+ N_VDD_X2/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X10/M7 N_X2/X10/9_X2/X10/M7_d N_X2/40_X2/X10/M7_g N_4_X2/X10/M7_s
+ N_VDD_X2/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X10/M8 N_VDD_X2/X10/M8_d N_X2/34_X2/X10/M8_g N_X2/X10/9_X2/X10/M8_s
+ N_VDD_X2/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X10/M9 N_VDD_X2/X10/M9_d N_4_X2/X10/M9_g N_46_X2/X10/M9_s N_VDD_X2/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X11/M0 N_GND_X2/X11/M0_d N_X2/X11/14_X2/X11/M0_g N_X2/X11/16_X2/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X11/M1 N_GND_X2/X11/M1_d N_X2/X11/13_X2/X11/M1_g N_X2/X11/14_X2/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X11/M2 N_X2/X11/20_X2/X11/M2_d N_B22_X2/X11/M2_g N_GND_X2/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X11/M3 N_X2/X11/14_X2/X11/M3_d N_A22_X2/X11/M3_g N_X2/X11/20_X2/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X11/M4 N_GND_X2/X11/M4_d N_X2/X11/13_X2/X11/M4_g N_X2/X11/17_X2/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X11/M5 N_X2/X11/13_X2/X11/M5_d N_B22_X2/X11/M5_g N_GND_X2/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X11/M6 N_GND_X2/X11/M6_d N_A22_X2/X11/M6_g N_X2/X11/13_X2/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X11/M7 N_X2/X11/15_X2/X11/M7_d N_X2/X11/13_X2/X11/M7_g
+ N_X2/X11/14_X2/X11/M7_s N_VDD_X2/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX2/X11/M8 N_VDD_X2/X11/M8_d N_B22_X2/X11/M8_g N_X2/X11/15_X2/X11/M8_s
+ N_VDD_X2/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X11/M9 N_X2/X11/15_X2/X11/M9_d N_A22_X2/X11/M9_g N_VDD_X2/X11/M9_s
+ N_VDD_X2/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X11/M10 N_VDD_X2/X11/M10_d N_X2/X11/14_X2/X11/M10_g N_X2/X11/16_X2/X11/M10_s
+ N_VDD_X2/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X11/M11 N_X2/X11/21_X2/X11/M11_d N_B22_X2/X11/M11_g N_VDD_X2/X11/M11_s
+ N_VDD_X2/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX2/X11/M12 N_X2/X11/13_X2/X11/M12_d N_A22_X2/X11/M12_g N_X2/X11/21_X2/X11/M12_s
+ N_VDD_X2/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X11/M13 N_VDD_X2/X11/M13_d N_X2/X11/13_X2/X11/M13_g N_X2/X11/17_X2/X11/M13_s
+ N_VDD_X2/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X11/X14/M0 N_GND_X2/X11/X14/M0_d N_X2/X11/18_X2/X11/X14/M0_g
+ N_SUM22_X2/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X11/X14/M1 N_X2/X11/X14/10_X2/X11/X14/M1_d N_X2/30_X2/X11/X14/M1_g
+ N_X2/X11/18_X2/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X11/X14/M2 N_GND_X2/X11/X14/M2_d N_X2/27_X2/X11/X14/M2_g
+ N_X2/X11/X14/10_X2/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X11/X14/M3 N_X2/X11/X14/11_X2/X11/X14/M3_d N_X2/X11/16_X2/X11/X14/M3_g
+ N_GND_X2/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X11/X14/M4 N_X2/X11/18_X2/X11/X14/M4_d N_X2/36_X2/X11/X14/M4_g
+ N_X2/X11/X14/11_X2/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X11/X14/M5 N_X2/X11/X14/9_X2/X11/X14/M5_d N_X2/X11/16_X2/X11/X14/M5_g
+ N_VDD_X2/X11/X14/M5_s N_VDD_X2/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X11/X14/M6 N_X2/X11/18_X2/X11/X14/M6_d N_X2/30_X2/X11/X14/M6_g
+ N_X2/X11/X14/9_X2/X11/X14/M6_s N_VDD_X2/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X14/M7 N_X2/X11/X14/9_X2/X11/X14/M7_d N_X2/27_X2/X11/X14/M7_g
+ N_X2/X11/18_X2/X11/X14/M7_s N_VDD_X2/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X14/M8 N_VDD_X2/X11/X14/M8_d N_X2/36_X2/X11/X14/M8_g
+ N_X2/X11/X14/9_X2/X11/X14/M8_s N_VDD_X2/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X11/X14/M9 N_VDD_X2/X11/X14/M9_d N_X2/X11/18_X2/X11/X14/M9_g
+ N_SUM22_X2/X11/X14/M9_s N_VDD_X2/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X11/X15/M0 N_GND_X2/X11/X15/M0_d N_X2/29_X2/X11/X15/M0_g
+ N_X2/38_X2/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X11/X15/M1 N_X2/X11/X15/10_X2/X11/X15/M1_d N_X2/X11/17_X2/X11/X15/M1_g
+ N_X2/29_X2/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX2/X11/X15/M2 N_GND_X2/X11/X15/M2_d N_X2/36_X2/X11/X15/M2_g
+ N_X2/X11/X15/10_X2/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X11/X15/M3 N_X2/X11/X15/11_X2/X11/X15/M3_d N_B22_X2/X11/X15/M3_g
+ N_GND_X2/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X11/X15/M4 N_X2/29_X2/X11/X15/M4_d N_A22_X2/X11/X15/M4_g
+ N_X2/X11/X15/11_X2/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X11/X15/M5 N_X2/X11/X15/9_X2/X11/X15/M5_d N_B22_X2/X11/X15/M5_g
+ N_VDD_X2/X11/X15/M5_s N_VDD_X2/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X11/X15/M6 N_X2/29_X2/X11/X15/M6_d N_X2/X11/17_X2/X11/X15/M6_g
+ N_X2/X11/X15/9_X2/X11/X15/M6_s N_VDD_X2/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X15/M7 N_X2/X11/X15/9_X2/X11/X15/M7_d N_X2/36_X2/X11/X15/M7_g
+ N_X2/29_X2/X11/X15/M7_s N_VDD_X2/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X15/M8 N_VDD_X2/X11/X15/M8_d N_A22_X2/X11/X15/M8_g
+ N_X2/X11/X15/9_X2/X11/X15/M8_s N_VDD_X2/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X11/X15/M9 N_VDD_X2/X11/X15/M9_d N_X2/29_X2/X11/X15/M9_g
+ N_X2/38_X2/X11/X15/M9_s N_VDD_X2/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X11/X16/M0 N_GND_X2/X11/X16/M0_d N_X2/X11/19_X2/X11/X16/M0_g
+ N_X2/30_X2/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X11/X16/M1 N_X2/X11/X16/10_X2/X11/X16/M1_d N_A22N_X2/X11/X16/M1_g
+ N_X2/X11/19_X2/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X11/X16/M2 N_GND_X2/X11/X16/M2_d N_B22_X2/X11/X16/M2_g
+ N_X2/X11/X16/10_X2/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X11/X16/M3 N_X2/X11/X16/11_X2/X11/X16/M3_d N_B22N_X2/X11/X16/M3_g
+ N_GND_X2/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X11/X16/M4 N_X2/X11/19_X2/X11/X16/M4_d N_A22_X2/X11/X16/M4_g
+ N_X2/X11/X16/11_X2/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X11/X16/M5 N_X2/X11/X16/9_X2/X11/X16/M5_d N_B22N_X2/X11/X16/M5_g
+ N_VDD_X2/X11/X16/M5_s N_VDD_X2/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X11/X16/M6 N_X2/X11/19_X2/X11/X16/M6_d N_A22N_X2/X11/X16/M6_g
+ N_X2/X11/X16/9_X2/X11/X16/M6_s N_VDD_X2/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X16/M7 N_X2/X11/X16/9_X2/X11/X16/M7_d N_B22_X2/X11/X16/M7_g
+ N_X2/X11/19_X2/X11/X16/M7_s N_VDD_X2/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X11/X16/M8 N_VDD_X2/X11/X16/M8_d N_A22_X2/X11/X16/M8_g
+ N_X2/X11/X16/9_X2/X11/X16/M8_s N_VDD_X2/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X11/X16/M9 N_VDD_X2/X11/X16/M9_d N_X2/X11/19_X2/X11/X16/M9_g
+ N_X2/30_X2/X11/X16/M9_s N_VDD_X2/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X12/M0 N_GND_X2/X12/M0_d N_X2/X12/14_X2/X12/M0_g N_X2/X12/16_X2/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X12/M1 N_GND_X2/X12/M1_d N_X2/X12/13_X2/X12/M1_g N_X2/X12/14_X2/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X12/M2 N_X2/X12/20_X2/X12/M2_d N_B21_X2/X12/M2_g N_GND_X2/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X12/M3 N_X2/X12/14_X2/X12/M3_d N_A21_X2/X12/M3_g N_X2/X12/20_X2/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X12/M4 N_GND_X2/X12/M4_d N_X2/X12/13_X2/X12/M4_g N_X2/X12/17_X2/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X12/M5 N_X2/X12/13_X2/X12/M5_d N_B21_X2/X12/M5_g N_GND_X2/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X12/M6 N_GND_X2/X12/M6_d N_A21_X2/X12/M6_g N_X2/X12/13_X2/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X12/M7 N_X2/X12/15_X2/X12/M7_d N_X2/X12/13_X2/X12/M7_g
+ N_X2/X12/14_X2/X12/M7_s N_VDD_X2/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX2/X12/M8 N_VDD_X2/X12/M8_d N_B21_X2/X12/M8_g N_X2/X12/15_X2/X12/M8_s
+ N_VDD_X2/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X12/M9 N_X2/X12/15_X2/X12/M9_d N_A21_X2/X12/M9_g N_VDD_X2/X12/M9_s
+ N_VDD_X2/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X12/M10 N_VDD_X2/X12/M10_d N_X2/X12/14_X2/X12/M10_g N_X2/X12/16_X2/X12/M10_s
+ N_VDD_X2/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X12/M11 N_X2/X12/21_X2/X12/M11_d N_B21_X2/X12/M11_g N_VDD_X2/X12/M11_s
+ N_VDD_X2/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX2/X12/M12 N_X2/X12/13_X2/X12/M12_d N_A21_X2/X12/M12_g N_X2/X12/21_X2/X12/M12_s
+ N_VDD_X2/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X12/M13 N_VDD_X2/X12/M13_d N_X2/X12/13_X2/X12/M13_g N_X2/X12/17_X2/X12/M13_s
+ N_VDD_X2/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X12/X14/M0 N_GND_X2/X12/X14/M0_d N_X2/X12/18_X2/X12/X14/M0_g
+ N_SUM21_X2/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X12/X14/M1 N_X2/X12/X14/10_X2/X12/X14/M1_d N_X2/31_X2/X12/X14/M1_g
+ N_X2/X12/18_X2/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X12/X14/M2 N_GND_X2/X12/X14/M2_d N_X2/28_X2/X12/X14/M2_g
+ N_X2/X12/X14/10_X2/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X12/X14/M3 N_X2/X12/X14/11_X2/X12/X14/M3_d N_X2/X12/16_X2/X12/X14/M3_g
+ N_GND_X2/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X12/X14/M4 N_X2/X12/18_X2/X12/X14/M4_d N_X2/37_X2/X12/X14/M4_g
+ N_X2/X12/X14/11_X2/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X12/X14/M5 N_X2/X12/X14/9_X2/X12/X14/M5_d N_X2/X12/16_X2/X12/X14/M5_g
+ N_VDD_X2/X12/X14/M5_s N_VDD_X2/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X12/X14/M6 N_X2/X12/18_X2/X12/X14/M6_d N_X2/31_X2/X12/X14/M6_g
+ N_X2/X12/X14/9_X2/X12/X14/M6_s N_VDD_X2/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X14/M7 N_X2/X12/X14/9_X2/X12/X14/M7_d N_X2/28_X2/X12/X14/M7_g
+ N_X2/X12/18_X2/X12/X14/M7_s N_VDD_X2/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X14/M8 N_VDD_X2/X12/X14/M8_d N_X2/37_X2/X12/X14/M8_g
+ N_X2/X12/X14/9_X2/X12/X14/M8_s N_VDD_X2/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X12/X14/M9 N_VDD_X2/X12/X14/M9_d N_X2/X12/18_X2/X12/X14/M9_g
+ N_SUM21_X2/X12/X14/M9_s N_VDD_X2/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X12/X15/M0 N_GND_X2/X12/X15/M0_d N_X2/27_X2/X12/X15/M0_g
+ N_X2/36_X2/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X12/X15/M1 N_X2/X12/X15/10_X2/X12/X15/M1_d N_X2/X12/17_X2/X12/X15/M1_g
+ N_X2/27_X2/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX2/X12/X15/M2 N_GND_X2/X12/X15/M2_d N_X2/37_X2/X12/X15/M2_g
+ N_X2/X12/X15/10_X2/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X12/X15/M3 N_X2/X12/X15/11_X2/X12/X15/M3_d N_B21_X2/X12/X15/M3_g
+ N_GND_X2/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X12/X15/M4 N_X2/27_X2/X12/X15/M4_d N_A21_X2/X12/X15/M4_g
+ N_X2/X12/X15/11_X2/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X12/X15/M5 N_X2/X12/X15/9_X2/X12/X15/M5_d N_B21_X2/X12/X15/M5_g
+ N_VDD_X2/X12/X15/M5_s N_VDD_X2/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X12/X15/M6 N_X2/27_X2/X12/X15/M6_d N_X2/X12/17_X2/X12/X15/M6_g
+ N_X2/X12/X15/9_X2/X12/X15/M6_s N_VDD_X2/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X15/M7 N_X2/X12/X15/9_X2/X12/X15/M7_d N_X2/37_X2/X12/X15/M7_g
+ N_X2/27_X2/X12/X15/M7_s N_VDD_X2/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X15/M8 N_VDD_X2/X12/X15/M8_d N_A21_X2/X12/X15/M8_g
+ N_X2/X12/X15/9_X2/X12/X15/M8_s N_VDD_X2/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X12/X15/M9 N_VDD_X2/X12/X15/M9_d N_X2/27_X2/X12/X15/M9_g
+ N_X2/36_X2/X12/X15/M9_s N_VDD_X2/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X12/X16/M0 N_GND_X2/X12/X16/M0_d N_X2/X12/19_X2/X12/X16/M0_g
+ N_X2/31_X2/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X12/X16/M1 N_X2/X12/X16/10_X2/X12/X16/M1_d N_A21N_X2/X12/X16/M1_g
+ N_X2/X12/19_X2/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X12/X16/M2 N_GND_X2/X12/X16/M2_d N_B21_X2/X12/X16/M2_g
+ N_X2/X12/X16/10_X2/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X12/X16/M3 N_X2/X12/X16/11_X2/X12/X16/M3_d N_B21N_X2/X12/X16/M3_g
+ N_GND_X2/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X12/X16/M4 N_X2/X12/19_X2/X12/X16/M4_d N_A21_X2/X12/X16/M4_g
+ N_X2/X12/X16/11_X2/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X12/X16/M5 N_X2/X12/X16/9_X2/X12/X16/M5_d N_B21N_X2/X12/X16/M5_g
+ N_VDD_X2/X12/X16/M5_s N_VDD_X2/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X12/X16/M6 N_X2/X12/19_X2/X12/X16/M6_d N_A21N_X2/X12/X16/M6_g
+ N_X2/X12/X16/9_X2/X12/X16/M6_s N_VDD_X2/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X16/M7 N_X2/X12/X16/9_X2/X12/X16/M7_d N_B21_X2/X12/X16/M7_g
+ N_X2/X12/19_X2/X12/X16/M7_s N_VDD_X2/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X12/X16/M8 N_VDD_X2/X12/X16/M8_d N_A21_X2/X12/X16/M8_g
+ N_X2/X12/X16/9_X2/X12/X16/M8_s N_VDD_X2/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X12/X16/M9 N_VDD_X2/X12/X16/M9_d N_X2/X12/19_X2/X12/X16/M9_g
+ N_X2/31_X2/X12/X16/M9_s N_VDD_X2/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X13/M0 N_GND_X2/X13/M0_d N_X2/X13/14_X2/X13/M0_g N_X2/X13/16_X2/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X13/M1 N_GND_X2/X13/M1_d N_X2/X13/13_X2/X13/M1_g N_X2/X13/14_X2/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X13/M2 N_X2/X13/20_X2/X13/M2_d N_B20_X2/X13/M2_g N_GND_X2/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X13/M3 N_X2/X13/14_X2/X13/M3_d N_A20_X2/X13/M3_g N_X2/X13/20_X2/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X13/M4 N_GND_X2/X13/M4_d N_X2/X13/13_X2/X13/M4_g N_X2/X13/17_X2/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X13/M5 N_X2/X13/13_X2/X13/M5_d N_B20_X2/X13/M5_g N_GND_X2/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X13/M6 N_GND_X2/X13/M6_d N_A20_X2/X13/M6_g N_X2/X13/13_X2/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X13/M7 N_X2/X13/15_X2/X13/M7_d N_X2/X13/13_X2/X13/M7_g
+ N_X2/X13/14_X2/X13/M7_s N_VDD_X2/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX2/X13/M8 N_VDD_X2/X13/M8_d N_B20_X2/X13/M8_g N_X2/X13/15_X2/X13/M8_s
+ N_VDD_X2/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X13/M9 N_X2/X13/15_X2/X13/M9_d N_A20_X2/X13/M9_g N_VDD_X2/X13/M9_s
+ N_VDD_X2/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X13/M10 N_VDD_X2/X13/M10_d N_X2/X13/14_X2/X13/M10_g N_X2/X13/16_X2/X13/M10_s
+ N_VDD_X2/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X13/M11 N_X2/X13/21_X2/X13/M11_d N_B20_X2/X13/M11_g N_VDD_X2/X13/M11_s
+ N_VDD_X2/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX2/X13/M12 N_X2/X13/13_X2/X13/M12_d N_A20_X2/X13/M12_g N_X2/X13/21_X2/X13/M12_s
+ N_VDD_X2/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X13/M13 N_VDD_X2/X13/M13_d N_X2/X13/13_X2/X13/M13_g N_X2/X13/17_X2/X13/M13_s
+ N_VDD_X2/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X13/X14/M0 N_GND_X2/X13/X14/M0_d N_X2/X13/18_X2/X13/X14/M0_g
+ N_SUM20_X2/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X13/X14/M1 N_X2/X13/X14/10_X2/X13/X14/M1_d N_X2/32_X2/X13/X14/M1_g
+ N_X2/X13/18_X2/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X13/X14/M2 N_GND_X2/X13/X14/M2_d N_5_X2/X13/X14/M2_g
+ N_X2/X13/X14/10_X2/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X13/X14/M3 N_X2/X13/X14/11_X2/X13/X14/M3_d N_X2/X13/16_X2/X13/X14/M3_g
+ N_GND_X2/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X13/X14/M4 N_X2/X13/18_X2/X13/X14/M4_d N_47_X2/X13/X14/M4_g
+ N_X2/X13/X14/11_X2/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X13/X14/M5 N_X2/X13/X14/9_X2/X13/X14/M5_d N_X2/X13/16_X2/X13/X14/M5_g
+ N_VDD_X2/X13/X14/M5_s N_VDD_X2/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X13/X14/M6 N_X2/X13/18_X2/X13/X14/M6_d N_X2/32_X2/X13/X14/M6_g
+ N_X2/X13/X14/9_X2/X13/X14/M6_s N_VDD_X2/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X14/M7 N_X2/X13/X14/9_X2/X13/X14/M7_d N_5_X2/X13/X14/M7_g
+ N_X2/X13/18_X2/X13/X14/M7_s N_VDD_X2/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X14/M8 N_VDD_X2/X13/X14/M8_d N_47_X2/X13/X14/M8_g
+ N_X2/X13/X14/9_X2/X13/X14/M8_s N_VDD_X2/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X13/X14/M9 N_VDD_X2/X13/X14/M9_d N_X2/X13/18_X2/X13/X14/M9_g
+ N_SUM20_X2/X13/X14/M9_s N_VDD_X2/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X13/X15/M0 N_GND_X2/X13/X15/M0_d N_X2/28_X2/X13/X15/M0_g
+ N_X2/37_X2/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X13/X15/M1 N_X2/X13/X15/10_X2/X13/X15/M1_d N_X2/X13/17_X2/X13/X15/M1_g
+ N_X2/28_X2/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX2/X13/X15/M2 N_GND_X2/X13/X15/M2_d N_47_X2/X13/X15/M2_g
+ N_X2/X13/X15/10_X2/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X13/X15/M3 N_X2/X13/X15/11_X2/X13/X15/M3_d N_B20_X2/X13/X15/M3_g
+ N_GND_X2/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X13/X15/M4 N_X2/28_X2/X13/X15/M4_d N_A20_X2/X13/X15/M4_g
+ N_X2/X13/X15/11_X2/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X13/X15/M5 N_X2/X13/X15/9_X2/X13/X15/M5_d N_B20_X2/X13/X15/M5_g
+ N_VDD_X2/X13/X15/M5_s N_VDD_X2/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X13/X15/M6 N_X2/28_X2/X13/X15/M6_d N_X2/X13/17_X2/X13/X15/M6_g
+ N_X2/X13/X15/9_X2/X13/X15/M6_s N_VDD_X2/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X15/M7 N_X2/X13/X15/9_X2/X13/X15/M7_d N_47_X2/X13/X15/M7_g
+ N_X2/28_X2/X13/X15/M7_s N_VDD_X2/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X15/M8 N_VDD_X2/X13/X15/M8_d N_A20_X2/X13/X15/M8_g
+ N_X2/X13/X15/9_X2/X13/X15/M8_s N_VDD_X2/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X13/X15/M9 N_VDD_X2/X13/X15/M9_d N_X2/28_X2/X13/X15/M9_g
+ N_X2/37_X2/X13/X15/M9_s N_VDD_X2/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X13/X16/M0 N_GND_X2/X13/X16/M0_d N_X2/X13/19_X2/X13/X16/M0_g
+ N_X2/32_X2/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X13/X16/M1 N_X2/X13/X16/10_X2/X13/X16/M1_d N_A20N_X2/X13/X16/M1_g
+ N_X2/X13/19_X2/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X13/X16/M2 N_GND_X2/X13/X16/M2_d N_B20_X2/X13/X16/M2_g
+ N_X2/X13/X16/10_X2/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X13/X16/M3 N_X2/X13/X16/11_X2/X13/X16/M3_d N_B20N_X2/X13/X16/M3_g
+ N_GND_X2/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X13/X16/M4 N_X2/X13/19_X2/X13/X16/M4_d N_A20_X2/X13/X16/M4_g
+ N_X2/X13/X16/11_X2/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X13/X16/M5 N_X2/X13/X16/9_X2/X13/X16/M5_d N_B20N_X2/X13/X16/M5_g
+ N_VDD_X2/X13/X16/M5_s N_VDD_X2/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X13/X16/M6 N_X2/X13/19_X2/X13/X16/M6_d N_A20N_X2/X13/X16/M6_g
+ N_X2/X13/X16/9_X2/X13/X16/M6_s N_VDD_X2/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X16/M7 N_X2/X13/X16/9_X2/X13/X16/M7_d N_B20_X2/X13/X16/M7_g
+ N_X2/X13/19_X2/X13/X16/M7_s N_VDD_X2/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X13/X16/M8 N_VDD_X2/X13/X16/M8_d N_A20_X2/X13/X16/M8_g
+ N_X2/X13/X16/9_X2/X13/X16/M8_s N_VDD_X2/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X13/X16/M9 N_VDD_X2/X13/X16/M9_d N_X2/X13/19_X2/X13/X16/M9_g
+ N_X2/32_X2/X13/X16/M9_s N_VDD_X2/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X14/M0 N_GND_X2/X14/M0_d N_X2/X14/14_X2/X14/M0_g N_X2/X14/16_X2/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X14/M1 N_GND_X2/X14/M1_d N_X2/X14/13_X2/X14/M1_g N_X2/X14/14_X2/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X14/M2 N_X2/X14/20_X2/X14/M2_d N_B23_X2/X14/M2_g N_GND_X2/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX2/X14/M3 N_X2/X14/14_X2/X14/M3_d N_A23_X2/X14/M3_g N_X2/X14/20_X2/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X14/M4 N_GND_X2/X14/M4_d N_X2/X14/13_X2/X14/M4_g N_X2/X14/17_X2/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X14/M5 N_X2/X14/13_X2/X14/M5_d N_B23_X2/X14/M5_g N_GND_X2/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX2/X14/M6 N_GND_X2/X14/M6_d N_A23_X2/X14/M6_g N_X2/X14/13_X2/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX2/X14/M7 N_X2/X14/15_X2/X14/M7_d N_X2/X14/13_X2/X14/M7_g
+ N_X2/X14/14_X2/X14/M7_s N_VDD_X2/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX2/X14/M8 N_VDD_X2/X14/M8_d N_B23_X2/X14/M8_g N_X2/X14/15_X2/X14/M8_s
+ N_VDD_X2/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX2/X14/M9 N_X2/X14/15_X2/X14/M9_d N_A23_X2/X14/M9_g N_VDD_X2/X14/M9_s
+ N_VDD_X2/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X14/M10 N_VDD_X2/X14/M10_d N_X2/X14/14_X2/X14/M10_g N_X2/X14/16_X2/X14/M10_s
+ N_VDD_X2/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X14/M11 N_X2/X14/21_X2/X14/M11_d N_B23_X2/X14/M11_g N_VDD_X2/X14/M11_s
+ N_VDD_X2/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX2/X14/M12 N_X2/X14/13_X2/X14/M12_d N_A23_X2/X14/M12_g N_X2/X14/21_X2/X14/M12_s
+ N_VDD_X2/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX2/X14/M13 N_VDD_X2/X14/M13_d N_X2/X14/13_X2/X14/M13_g N_X2/X14/17_X2/X14/M13_s
+ N_VDD_X2/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X14/X14/M0 N_GND_X2/X14/X14/M0_d N_X2/X14/18_X2/X14/X14/M0_g
+ N_SUM23_X2/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X14/X14/M1 N_X2/X14/X14/10_X2/X14/X14/M1_d N_X2/35_X2/X14/X14/M1_g
+ N_X2/X14/18_X2/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X14/X14/M2 N_GND_X2/X14/X14/M2_d N_X2/29_X2/X14/X14/M2_g
+ N_X2/X14/X14/10_X2/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X14/X14/M3 N_X2/X14/X14/11_X2/X14/X14/M3_d N_X2/X14/16_X2/X14/X14/M3_g
+ N_GND_X2/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X14/X14/M4 N_X2/X14/18_X2/X14/X14/M4_d N_X2/38_X2/X14/X14/M4_g
+ N_X2/X14/X14/11_X2/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X14/X14/M5 N_X2/X14/X14/9_X2/X14/X14/M5_d N_X2/X14/16_X2/X14/X14/M5_g
+ N_VDD_X2/X14/X14/M5_s N_VDD_X2/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X14/X14/M6 N_X2/X14/18_X2/X14/X14/M6_d N_X2/35_X2/X14/X14/M6_g
+ N_X2/X14/X14/9_X2/X14/X14/M6_s N_VDD_X2/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X14/M7 N_X2/X14/X14/9_X2/X14/X14/M7_d N_X2/29_X2/X14/X14/M7_g
+ N_X2/X14/18_X2/X14/X14/M7_s N_VDD_X2/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X14/M8 N_VDD_X2/X14/X14/M8_d N_X2/38_X2/X14/X14/M8_g
+ N_X2/X14/X14/9_X2/X14/X14/M8_s N_VDD_X2/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X14/X14/M9 N_VDD_X2/X14/X14/M9_d N_X2/X14/18_X2/X14/X14/M9_g
+ N_SUM23_X2/X14/X14/M9_s N_VDD_X2/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X14/X15/M0 N_GND_X2/X14/X15/M0_d N_X2/33_X2/X14/X15/M0_g
+ N_X2/34_X2/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X14/X15/M1 N_X2/X14/X15/10_X2/X14/X15/M1_d N_X2/X14/17_X2/X14/X15/M1_g
+ N_X2/33_X2/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX2/X14/X15/M2 N_GND_X2/X14/X15/M2_d N_X2/38_X2/X14/X15/M2_g
+ N_X2/X14/X15/10_X2/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X14/X15/M3 N_X2/X14/X15/11_X2/X14/X15/M3_d N_B23_X2/X14/X15/M3_g
+ N_GND_X2/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X14/X15/M4 N_X2/33_X2/X14/X15/M4_d N_A23_X2/X14/X15/M4_g
+ N_X2/X14/X15/11_X2/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X14/X15/M5 N_X2/X14/X15/9_X2/X14/X15/M5_d N_B23_X2/X14/X15/M5_g
+ N_VDD_X2/X14/X15/M5_s N_VDD_X2/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X14/X15/M6 N_X2/33_X2/X14/X15/M6_d N_X2/X14/17_X2/X14/X15/M6_g
+ N_X2/X14/X15/9_X2/X14/X15/M6_s N_VDD_X2/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X15/M7 N_X2/X14/X15/9_X2/X14/X15/M7_d N_X2/38_X2/X14/X15/M7_g
+ N_X2/33_X2/X14/X15/M7_s N_VDD_X2/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X15/M8 N_VDD_X2/X14/X15/M8_d N_A23_X2/X14/X15/M8_g
+ N_X2/X14/X15/9_X2/X14/X15/M8_s N_VDD_X2/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X14/X15/M9 N_VDD_X2/X14/X15/M9_d N_X2/33_X2/X14/X15/M9_g
+ N_X2/34_X2/X14/X15/M9_s N_VDD_X2/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX2/X14/X16/M0 N_GND_X2/X14/X16/M0_d N_X2/X14/19_X2/X14/X16/M0_g
+ N_X2/35_X2/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX2/X14/X16/M1 N_X2/X14/X16/10_X2/X14/X16/M1_d N_A23N_X2/X14/X16/M1_g
+ N_X2/X14/19_X2/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX2/X14/X16/M2 N_GND_X2/X14/X16/M2_d N_B23_X2/X14/X16/M2_g
+ N_X2/X14/X16/10_X2/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX2/X14/X16/M3 N_X2/X14/X16/11_X2/X14/X16/M3_d N_B23N_X2/X14/X16/M3_g
+ N_GND_X2/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX2/X14/X16/M4 N_X2/X14/19_X2/X14/X16/M4_d N_A23_X2/X14/X16/M4_g
+ N_X2/X14/X16/11_X2/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX2/X14/X16/M5 N_X2/X14/X16/9_X2/X14/X16/M5_d N_B23N_X2/X14/X16/M5_g
+ N_VDD_X2/X14/X16/M5_s N_VDD_X2/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX2/X14/X16/M6 N_X2/X14/19_X2/X14/X16/M6_d N_A23N_X2/X14/X16/M6_g
+ N_X2/X14/X16/9_X2/X14/X16/M6_s N_VDD_X2/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X16/M7 N_X2/X14/X16/9_X2/X14/X16/M7_d N_B23_X2/X14/X16/M7_g
+ N_X2/X14/19_X2/X14/X16/M7_s N_VDD_X2/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX2/X14/X16/M8 N_VDD_X2/X14/X16/M8_d N_A23_X2/X14/X16/M8_g
+ N_X2/X14/X16/9_X2/X14/X16/M8_s N_VDD_X2/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX2/X14/X16/M9 N_VDD_X2/X14/X16/M9_d N_X2/X14/19_X2/X14/X16/M9_g
+ N_X2/35_X2/X14/X16/M9_s N_VDD_X2/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/M0 N_GND_X3/M0_d N_X3/39_X3/M0_g N_X3/40_X3/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/M1 N_X3/41_X3/M1_d N_X3/32_X3/M1_g N_GND_X3/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX3/M2 N_X3/42_X3/M2_d N_X3/31_X3/M2_g N_X3/41_X3/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX3/M3 N_X3/43_X3/M3_d N_X3/30_X3/M3_g N_X3/42_X3/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX3/M4 N_X3/39_X3/M4_d N_X3/35_X3/M4_g N_X3/43_X3/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX3/M5 N_VDD_X3/M5_d N_X3/39_X3/M5_g N_X3/40_X3/M5_s N_VDD_X3/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/M6 N_X3/39_X3/M6_d N_X3/32_X3/M6_g N_VDD_X3/M6_s N_VDD_X3/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX3/M7 N_VDD_X3/M7_d N_X3/31_X3/M7_g N_X3/39_X3/M7_s N_VDD_X3/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX3/M8 N_X3/39_X3/M8_d N_X3/30_X3/M8_g N_VDD_X3/M8_s N_VDD_X3/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX3/M9 N_VDD_X3/M9_d N_X3/35_X3/M9_g N_X3/39_X3/M9_s N_VDD_X3/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX3/X10/M0 N_GND_X3/X10/M0_d N_8_X3/X10/M0_g N_50_X3/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X10/M1 N_X3/X10/10_X3/X10/M1_d N_48_X3/X10/M1_g N_8_X3/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X10/M2 N_GND_X3/X10/M2_d N_X3/40_X3/X10/M2_g N_X3/X10/10_X3/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X10/M3 N_X3/X10/11_X3/X10/M3_d N_X3/39_X3/X10/M3_g N_GND_X3/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X10/M4 N_8_X3/X10/M4_d N_X3/34_X3/X10/M4_g N_X3/X10/11_X3/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X10/M5 N_X3/X10/9_X3/X10/M5_d N_X3/39_X3/X10/M5_g N_VDD_X3/X10/M5_s
+ N_VDD_X3/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX3/X10/M6 N_8_X3/X10/M6_d N_48_X3/X10/M6_g N_X3/X10/9_X3/X10/M6_s
+ N_VDD_X3/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X10/M7 N_X3/X10/9_X3/X10/M7_d N_X3/40_X3/X10/M7_g N_8_X3/X10/M7_s
+ N_VDD_X3/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X10/M8 N_VDD_X3/X10/M8_d N_X3/34_X3/X10/M8_g N_X3/X10/9_X3/X10/M8_s
+ N_VDD_X3/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X10/M9 N_VDD_X3/X10/M9_d N_8_X3/X10/M9_g N_50_X3/X10/M9_s N_VDD_X3/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X11/M0 N_GND_X3/X11/M0_d N_X3/X11/14_X3/X11/M0_g N_X3/X11/16_X3/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X11/M1 N_GND_X3/X11/M1_d N_X3/X11/13_X3/X11/M1_g N_X3/X11/14_X3/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X11/M2 N_X3/X11/20_X3/X11/M2_d N_B14_X3/X11/M2_g N_GND_X3/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X11/M3 N_X3/X11/14_X3/X11/M3_d N_A14_X3/X11/M3_g N_X3/X11/20_X3/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X11/M4 N_GND_X3/X11/M4_d N_X3/X11/13_X3/X11/M4_g N_X3/X11/17_X3/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X11/M5 N_X3/X11/13_X3/X11/M5_d N_B14_X3/X11/M5_g N_GND_X3/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X11/M6 N_GND_X3/X11/M6_d N_A14_X3/X11/M6_g N_X3/X11/13_X3/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X11/M7 N_X3/X11/15_X3/X11/M7_d N_X3/X11/13_X3/X11/M7_g
+ N_X3/X11/14_X3/X11/M7_s N_VDD_X3/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX3/X11/M8 N_VDD_X3/X11/M8_d N_B14_X3/X11/M8_g N_X3/X11/15_X3/X11/M8_s
+ N_VDD_X3/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X11/M9 N_X3/X11/15_X3/X11/M9_d N_A14_X3/X11/M9_g N_VDD_X3/X11/M9_s
+ N_VDD_X3/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X11/M10 N_VDD_X3/X11/M10_d N_X3/X11/14_X3/X11/M10_g N_X3/X11/16_X3/X11/M10_s
+ N_VDD_X3/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X11/M11 N_X3/X11/21_X3/X11/M11_d N_B14_X3/X11/M11_g N_VDD_X3/X11/M11_s
+ N_VDD_X3/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX3/X11/M12 N_X3/X11/13_X3/X11/M12_d N_A14_X3/X11/M12_g N_X3/X11/21_X3/X11/M12_s
+ N_VDD_X3/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X11/M13 N_VDD_X3/X11/M13_d N_X3/X11/13_X3/X11/M13_g N_X3/X11/17_X3/X11/M13_s
+ N_VDD_X3/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X11/X14/M0 N_GND_X3/X11/X14/M0_d N_X3/X11/18_X3/X11/X14/M0_g
+ N_SUM14_X3/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X11/X14/M1 N_X3/X11/X14/10_X3/X11/X14/M1_d N_X3/30_X3/X11/X14/M1_g
+ N_X3/X11/18_X3/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X11/X14/M2 N_GND_X3/X11/X14/M2_d N_X3/27_X3/X11/X14/M2_g
+ N_X3/X11/X14/10_X3/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X11/X14/M3 N_X3/X11/X14/11_X3/X11/X14/M3_d N_X3/X11/16_X3/X11/X14/M3_g
+ N_GND_X3/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X11/X14/M4 N_X3/X11/18_X3/X11/X14/M4_d N_X3/36_X3/X11/X14/M4_g
+ N_X3/X11/X14/11_X3/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X11/X14/M5 N_X3/X11/X14/9_X3/X11/X14/M5_d N_X3/X11/16_X3/X11/X14/M5_g
+ N_VDD_X3/X11/X14/M5_s N_VDD_X3/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X11/X14/M6 N_X3/X11/18_X3/X11/X14/M6_d N_X3/30_X3/X11/X14/M6_g
+ N_X3/X11/X14/9_X3/X11/X14/M6_s N_VDD_X3/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X14/M7 N_X3/X11/X14/9_X3/X11/X14/M7_d N_X3/27_X3/X11/X14/M7_g
+ N_X3/X11/18_X3/X11/X14/M7_s N_VDD_X3/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X14/M8 N_VDD_X3/X11/X14/M8_d N_X3/36_X3/X11/X14/M8_g
+ N_X3/X11/X14/9_X3/X11/X14/M8_s N_VDD_X3/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X11/X14/M9 N_VDD_X3/X11/X14/M9_d N_X3/X11/18_X3/X11/X14/M9_g
+ N_SUM14_X3/X11/X14/M9_s N_VDD_X3/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X11/X15/M0 N_GND_X3/X11/X15/M0_d N_X3/29_X3/X11/X15/M0_g
+ N_X3/38_X3/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X11/X15/M1 N_X3/X11/X15/10_X3/X11/X15/M1_d N_X3/X11/17_X3/X11/X15/M1_g
+ N_X3/29_X3/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX3/X11/X15/M2 N_GND_X3/X11/X15/M2_d N_X3/36_X3/X11/X15/M2_g
+ N_X3/X11/X15/10_X3/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X11/X15/M3 N_X3/X11/X15/11_X3/X11/X15/M3_d N_B14_X3/X11/X15/M3_g
+ N_GND_X3/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X11/X15/M4 N_X3/29_X3/X11/X15/M4_d N_A14_X3/X11/X15/M4_g
+ N_X3/X11/X15/11_X3/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X11/X15/M5 N_X3/X11/X15/9_X3/X11/X15/M5_d N_B14_X3/X11/X15/M5_g
+ N_VDD_X3/X11/X15/M5_s N_VDD_X3/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X11/X15/M6 N_X3/29_X3/X11/X15/M6_d N_X3/X11/17_X3/X11/X15/M6_g
+ N_X3/X11/X15/9_X3/X11/X15/M6_s N_VDD_X3/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X15/M7 N_X3/X11/X15/9_X3/X11/X15/M7_d N_X3/36_X3/X11/X15/M7_g
+ N_X3/29_X3/X11/X15/M7_s N_VDD_X3/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X15/M8 N_VDD_X3/X11/X15/M8_d N_A14_X3/X11/X15/M8_g
+ N_X3/X11/X15/9_X3/X11/X15/M8_s N_VDD_X3/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X11/X15/M9 N_VDD_X3/X11/X15/M9_d N_X3/29_X3/X11/X15/M9_g
+ N_X3/38_X3/X11/X15/M9_s N_VDD_X3/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X11/X16/M0 N_GND_X3/X11/X16/M0_d N_X3/X11/19_X3/X11/X16/M0_g
+ N_X3/30_X3/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X11/X16/M1 N_X3/X11/X16/10_X3/X11/X16/M1_d N_A14N_X3/X11/X16/M1_g
+ N_X3/X11/19_X3/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X11/X16/M2 N_GND_X3/X11/X16/M2_d N_B14_X3/X11/X16/M2_g
+ N_X3/X11/X16/10_X3/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X11/X16/M3 N_X3/X11/X16/11_X3/X11/X16/M3_d N_B14N_X3/X11/X16/M3_g
+ N_GND_X3/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X11/X16/M4 N_X3/X11/19_X3/X11/X16/M4_d N_A14_X3/X11/X16/M4_g
+ N_X3/X11/X16/11_X3/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X11/X16/M5 N_X3/X11/X16/9_X3/X11/X16/M5_d N_B14N_X3/X11/X16/M5_g
+ N_VDD_X3/X11/X16/M5_s N_VDD_X3/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X11/X16/M6 N_X3/X11/19_X3/X11/X16/M6_d N_A14N_X3/X11/X16/M6_g
+ N_X3/X11/X16/9_X3/X11/X16/M6_s N_VDD_X3/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X16/M7 N_X3/X11/X16/9_X3/X11/X16/M7_d N_B14_X3/X11/X16/M7_g
+ N_X3/X11/19_X3/X11/X16/M7_s N_VDD_X3/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X11/X16/M8 N_VDD_X3/X11/X16/M8_d N_A14_X3/X11/X16/M8_g
+ N_X3/X11/X16/9_X3/X11/X16/M8_s N_VDD_X3/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X11/X16/M9 N_VDD_X3/X11/X16/M9_d N_X3/X11/19_X3/X11/X16/M9_g
+ N_X3/30_X3/X11/X16/M9_s N_VDD_X3/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X12/M0 N_GND_X3/X12/M0_d N_X3/X12/14_X3/X12/M0_g N_X3/X12/16_X3/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X12/M1 N_GND_X3/X12/M1_d N_X3/X12/13_X3/X12/M1_g N_X3/X12/14_X3/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X12/M2 N_X3/X12/20_X3/X12/M2_d N_B13_X3/X12/M2_g N_GND_X3/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X12/M3 N_X3/X12/14_X3/X12/M3_d N_A13_X3/X12/M3_g N_X3/X12/20_X3/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X12/M4 N_GND_X3/X12/M4_d N_X3/X12/13_X3/X12/M4_g N_X3/X12/17_X3/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X12/M5 N_X3/X12/13_X3/X12/M5_d N_B13_X3/X12/M5_g N_GND_X3/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X12/M6 N_GND_X3/X12/M6_d N_A13_X3/X12/M6_g N_X3/X12/13_X3/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X12/M7 N_X3/X12/15_X3/X12/M7_d N_X3/X12/13_X3/X12/M7_g
+ N_X3/X12/14_X3/X12/M7_s N_VDD_X3/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX3/X12/M8 N_VDD_X3/X12/M8_d N_B13_X3/X12/M8_g N_X3/X12/15_X3/X12/M8_s
+ N_VDD_X3/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X12/M9 N_X3/X12/15_X3/X12/M9_d N_A13_X3/X12/M9_g N_VDD_X3/X12/M9_s
+ N_VDD_X3/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X12/M10 N_VDD_X3/X12/M10_d N_X3/X12/14_X3/X12/M10_g N_X3/X12/16_X3/X12/M10_s
+ N_VDD_X3/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X12/M11 N_X3/X12/21_X3/X12/M11_d N_B13_X3/X12/M11_g N_VDD_X3/X12/M11_s
+ N_VDD_X3/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX3/X12/M12 N_X3/X12/13_X3/X12/M12_d N_A13_X3/X12/M12_g N_X3/X12/21_X3/X12/M12_s
+ N_VDD_X3/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X12/M13 N_VDD_X3/X12/M13_d N_X3/X12/13_X3/X12/M13_g N_X3/X12/17_X3/X12/M13_s
+ N_VDD_X3/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X12/X14/M0 N_GND_X3/X12/X14/M0_d N_X3/X12/18_X3/X12/X14/M0_g
+ N_SUM13_X3/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X12/X14/M1 N_X3/X12/X14/10_X3/X12/X14/M1_d N_X3/31_X3/X12/X14/M1_g
+ N_X3/X12/18_X3/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X12/X14/M2 N_GND_X3/X12/X14/M2_d N_X3/28_X3/X12/X14/M2_g
+ N_X3/X12/X14/10_X3/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X12/X14/M3 N_X3/X12/X14/11_X3/X12/X14/M3_d N_X3/X12/16_X3/X12/X14/M3_g
+ N_GND_X3/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X12/X14/M4 N_X3/X12/18_X3/X12/X14/M4_d N_X3/37_X3/X12/X14/M4_g
+ N_X3/X12/X14/11_X3/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X12/X14/M5 N_X3/X12/X14/9_X3/X12/X14/M5_d N_X3/X12/16_X3/X12/X14/M5_g
+ N_VDD_X3/X12/X14/M5_s N_VDD_X3/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X12/X14/M6 N_X3/X12/18_X3/X12/X14/M6_d N_X3/31_X3/X12/X14/M6_g
+ N_X3/X12/X14/9_X3/X12/X14/M6_s N_VDD_X3/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X14/M7 N_X3/X12/X14/9_X3/X12/X14/M7_d N_X3/28_X3/X12/X14/M7_g
+ N_X3/X12/18_X3/X12/X14/M7_s N_VDD_X3/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X14/M8 N_VDD_X3/X12/X14/M8_d N_X3/37_X3/X12/X14/M8_g
+ N_X3/X12/X14/9_X3/X12/X14/M8_s N_VDD_X3/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X12/X14/M9 N_VDD_X3/X12/X14/M9_d N_X3/X12/18_X3/X12/X14/M9_g
+ N_SUM13_X3/X12/X14/M9_s N_VDD_X3/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X12/X15/M0 N_GND_X3/X12/X15/M0_d N_X3/27_X3/X12/X15/M0_g
+ N_X3/36_X3/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X12/X15/M1 N_X3/X12/X15/10_X3/X12/X15/M1_d N_X3/X12/17_X3/X12/X15/M1_g
+ N_X3/27_X3/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX3/X12/X15/M2 N_GND_X3/X12/X15/M2_d N_X3/37_X3/X12/X15/M2_g
+ N_X3/X12/X15/10_X3/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X12/X15/M3 N_X3/X12/X15/11_X3/X12/X15/M3_d N_B13_X3/X12/X15/M3_g
+ N_GND_X3/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X12/X15/M4 N_X3/27_X3/X12/X15/M4_d N_A13_X3/X12/X15/M4_g
+ N_X3/X12/X15/11_X3/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X12/X15/M5 N_X3/X12/X15/9_X3/X12/X15/M5_d N_B13_X3/X12/X15/M5_g
+ N_VDD_X3/X12/X15/M5_s N_VDD_X3/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X12/X15/M6 N_X3/27_X3/X12/X15/M6_d N_X3/X12/17_X3/X12/X15/M6_g
+ N_X3/X12/X15/9_X3/X12/X15/M6_s N_VDD_X3/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X15/M7 N_X3/X12/X15/9_X3/X12/X15/M7_d N_X3/37_X3/X12/X15/M7_g
+ N_X3/27_X3/X12/X15/M7_s N_VDD_X3/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X15/M8 N_VDD_X3/X12/X15/M8_d N_A13_X3/X12/X15/M8_g
+ N_X3/X12/X15/9_X3/X12/X15/M8_s N_VDD_X3/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X12/X15/M9 N_VDD_X3/X12/X15/M9_d N_X3/27_X3/X12/X15/M9_g
+ N_X3/36_X3/X12/X15/M9_s N_VDD_X3/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X12/X16/M0 N_GND_X3/X12/X16/M0_d N_X3/X12/19_X3/X12/X16/M0_g
+ N_X3/31_X3/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X12/X16/M1 N_X3/X12/X16/10_X3/X12/X16/M1_d N_A13N_X3/X12/X16/M1_g
+ N_X3/X12/19_X3/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X12/X16/M2 N_GND_X3/X12/X16/M2_d N_B13_X3/X12/X16/M2_g
+ N_X3/X12/X16/10_X3/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X12/X16/M3 N_X3/X12/X16/11_X3/X12/X16/M3_d N_B13N_X3/X12/X16/M3_g
+ N_GND_X3/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X12/X16/M4 N_X3/X12/19_X3/X12/X16/M4_d N_A13_X3/X12/X16/M4_g
+ N_X3/X12/X16/11_X3/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X12/X16/M5 N_X3/X12/X16/9_X3/X12/X16/M5_d N_B13N_X3/X12/X16/M5_g
+ N_VDD_X3/X12/X16/M5_s N_VDD_X3/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X12/X16/M6 N_X3/X12/19_X3/X12/X16/M6_d N_A13N_X3/X12/X16/M6_g
+ N_X3/X12/X16/9_X3/X12/X16/M6_s N_VDD_X3/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X16/M7 N_X3/X12/X16/9_X3/X12/X16/M7_d N_B13_X3/X12/X16/M7_g
+ N_X3/X12/19_X3/X12/X16/M7_s N_VDD_X3/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X12/X16/M8 N_VDD_X3/X12/X16/M8_d N_A13_X3/X12/X16/M8_g
+ N_X3/X12/X16/9_X3/X12/X16/M8_s N_VDD_X3/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X12/X16/M9 N_VDD_X3/X12/X16/M9_d N_X3/X12/19_X3/X12/X16/M9_g
+ N_X3/31_X3/X12/X16/M9_s N_VDD_X3/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X13/M0 N_GND_X3/X13/M0_d N_X3/X13/14_X3/X13/M0_g N_X3/X13/16_X3/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X13/M1 N_GND_X3/X13/M1_d N_X3/X13/13_X3/X13/M1_g N_X3/X13/14_X3/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X13/M2 N_X3/X13/20_X3/X13/M2_d N_B12_X3/X13/M2_g N_GND_X3/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X13/M3 N_X3/X13/14_X3/X13/M3_d N_A12_X3/X13/M3_g N_X3/X13/20_X3/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X13/M4 N_GND_X3/X13/M4_d N_X3/X13/13_X3/X13/M4_g N_X3/X13/17_X3/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X13/M5 N_X3/X13/13_X3/X13/M5_d N_B12_X3/X13/M5_g N_GND_X3/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X13/M6 N_GND_X3/X13/M6_d N_A12_X3/X13/M6_g N_X3/X13/13_X3/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X13/M7 N_X3/X13/15_X3/X13/M7_d N_X3/X13/13_X3/X13/M7_g
+ N_X3/X13/14_X3/X13/M7_s N_VDD_X3/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX3/X13/M8 N_VDD_X3/X13/M8_d N_B12_X3/X13/M8_g N_X3/X13/15_X3/X13/M8_s
+ N_VDD_X3/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X13/M9 N_X3/X13/15_X3/X13/M9_d N_A12_X3/X13/M9_g N_VDD_X3/X13/M9_s
+ N_VDD_X3/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X13/M10 N_VDD_X3/X13/M10_d N_X3/X13/14_X3/X13/M10_g N_X3/X13/16_X3/X13/M10_s
+ N_VDD_X3/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X13/M11 N_X3/X13/21_X3/X13/M11_d N_B12_X3/X13/M11_g N_VDD_X3/X13/M11_s
+ N_VDD_X3/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX3/X13/M12 N_X3/X13/13_X3/X13/M12_d N_A12_X3/X13/M12_g N_X3/X13/21_X3/X13/M12_s
+ N_VDD_X3/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X13/M13 N_VDD_X3/X13/M13_d N_X3/X13/13_X3/X13/M13_g N_X3/X13/17_X3/X13/M13_s
+ N_VDD_X3/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X13/X14/M0 N_GND_X3/X13/X14/M0_d N_X3/X13/18_X3/X13/X14/M0_g
+ N_SUM12_X3/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X13/X14/M1 N_X3/X13/X14/10_X3/X13/X14/M1_d N_X3/32_X3/X13/X14/M1_g
+ N_X3/X13/18_X3/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X13/X14/M2 N_GND_X3/X13/X14/M2_d N_6_X3/X13/X14/M2_g
+ N_X3/X13/X14/10_X3/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X13/X14/M3 N_X3/X13/X14/11_X3/X13/X14/M3_d N_X3/X13/16_X3/X13/X14/M3_g
+ N_GND_X3/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X13/X14/M4 N_X3/X13/18_X3/X13/X14/M4_d N_48_X3/X13/X14/M4_g
+ N_X3/X13/X14/11_X3/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X13/X14/M5 N_X3/X13/X14/9_X3/X13/X14/M5_d N_X3/X13/16_X3/X13/X14/M5_g
+ N_VDD_X3/X13/X14/M5_s N_VDD_X3/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X13/X14/M6 N_X3/X13/18_X3/X13/X14/M6_d N_X3/32_X3/X13/X14/M6_g
+ N_X3/X13/X14/9_X3/X13/X14/M6_s N_VDD_X3/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X14/M7 N_X3/X13/X14/9_X3/X13/X14/M7_d N_6_X3/X13/X14/M7_g
+ N_X3/X13/18_X3/X13/X14/M7_s N_VDD_X3/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X14/M8 N_VDD_X3/X13/X14/M8_d N_48_X3/X13/X14/M8_g
+ N_X3/X13/X14/9_X3/X13/X14/M8_s N_VDD_X3/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X13/X14/M9 N_VDD_X3/X13/X14/M9_d N_X3/X13/18_X3/X13/X14/M9_g
+ N_SUM12_X3/X13/X14/M9_s N_VDD_X3/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X13/X15/M0 N_GND_X3/X13/X15/M0_d N_X3/28_X3/X13/X15/M0_g
+ N_X3/37_X3/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X13/X15/M1 N_X3/X13/X15/10_X3/X13/X15/M1_d N_X3/X13/17_X3/X13/X15/M1_g
+ N_X3/28_X3/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX3/X13/X15/M2 N_GND_X3/X13/X15/M2_d N_48_X3/X13/X15/M2_g
+ N_X3/X13/X15/10_X3/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X13/X15/M3 N_X3/X13/X15/11_X3/X13/X15/M3_d N_B12_X3/X13/X15/M3_g
+ N_GND_X3/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X13/X15/M4 N_X3/28_X3/X13/X15/M4_d N_A12_X3/X13/X15/M4_g
+ N_X3/X13/X15/11_X3/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X13/X15/M5 N_X3/X13/X15/9_X3/X13/X15/M5_d N_B12_X3/X13/X15/M5_g
+ N_VDD_X3/X13/X15/M5_s N_VDD_X3/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X13/X15/M6 N_X3/28_X3/X13/X15/M6_d N_X3/X13/17_X3/X13/X15/M6_g
+ N_X3/X13/X15/9_X3/X13/X15/M6_s N_VDD_X3/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X15/M7 N_X3/X13/X15/9_X3/X13/X15/M7_d N_48_X3/X13/X15/M7_g
+ N_X3/28_X3/X13/X15/M7_s N_VDD_X3/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X15/M8 N_VDD_X3/X13/X15/M8_d N_A12_X3/X13/X15/M8_g
+ N_X3/X13/X15/9_X3/X13/X15/M8_s N_VDD_X3/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X13/X15/M9 N_VDD_X3/X13/X15/M9_d N_X3/28_X3/X13/X15/M9_g
+ N_X3/37_X3/X13/X15/M9_s N_VDD_X3/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X13/X16/M0 N_GND_X3/X13/X16/M0_d N_X3/X13/19_X3/X13/X16/M0_g
+ N_X3/32_X3/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X13/X16/M1 N_X3/X13/X16/10_X3/X13/X16/M1_d N_A12N_X3/X13/X16/M1_g
+ N_X3/X13/19_X3/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X13/X16/M2 N_GND_X3/X13/X16/M2_d N_B12_X3/X13/X16/M2_g
+ N_X3/X13/X16/10_X3/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X13/X16/M3 N_X3/X13/X16/11_X3/X13/X16/M3_d N_B12N_X3/X13/X16/M3_g
+ N_GND_X3/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X13/X16/M4 N_X3/X13/19_X3/X13/X16/M4_d N_A12_X3/X13/X16/M4_g
+ N_X3/X13/X16/11_X3/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X13/X16/M5 N_X3/X13/X16/9_X3/X13/X16/M5_d N_B12N_X3/X13/X16/M5_g
+ N_VDD_X3/X13/X16/M5_s N_VDD_X3/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X13/X16/M6 N_X3/X13/19_X3/X13/X16/M6_d N_A12N_X3/X13/X16/M6_g
+ N_X3/X13/X16/9_X3/X13/X16/M6_s N_VDD_X3/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X16/M7 N_X3/X13/X16/9_X3/X13/X16/M7_d N_B12_X3/X13/X16/M7_g
+ N_X3/X13/19_X3/X13/X16/M7_s N_VDD_X3/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X13/X16/M8 N_VDD_X3/X13/X16/M8_d N_A12_X3/X13/X16/M8_g
+ N_X3/X13/X16/9_X3/X13/X16/M8_s N_VDD_X3/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X13/X16/M9 N_VDD_X3/X13/X16/M9_d N_X3/X13/19_X3/X13/X16/M9_g
+ N_X3/32_X3/X13/X16/M9_s N_VDD_X3/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X14/M0 N_GND_X3/X14/M0_d N_X3/X14/14_X3/X14/M0_g N_X3/X14/16_X3/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X14/M1 N_GND_X3/X14/M1_d N_X3/X14/13_X3/X14/M1_g N_X3/X14/14_X3/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X14/M2 N_X3/X14/20_X3/X14/M2_d N_B15_X3/X14/M2_g N_GND_X3/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX3/X14/M3 N_X3/X14/14_X3/X14/M3_d N_A15_X3/X14/M3_g N_X3/X14/20_X3/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X14/M4 N_GND_X3/X14/M4_d N_X3/X14/13_X3/X14/M4_g N_X3/X14/17_X3/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X14/M5 N_X3/X14/13_X3/X14/M5_d N_B15_X3/X14/M5_g N_GND_X3/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX3/X14/M6 N_GND_X3/X14/M6_d N_A15_X3/X14/M6_g N_X3/X14/13_X3/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX3/X14/M7 N_X3/X14/15_X3/X14/M7_d N_X3/X14/13_X3/X14/M7_g
+ N_X3/X14/14_X3/X14/M7_s N_VDD_X3/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX3/X14/M8 N_VDD_X3/X14/M8_d N_B15_X3/X14/M8_g N_X3/X14/15_X3/X14/M8_s
+ N_VDD_X3/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX3/X14/M9 N_X3/X14/15_X3/X14/M9_d N_A15_X3/X14/M9_g N_VDD_X3/X14/M9_s
+ N_VDD_X3/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X14/M10 N_VDD_X3/X14/M10_d N_X3/X14/14_X3/X14/M10_g N_X3/X14/16_X3/X14/M10_s
+ N_VDD_X3/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X14/M11 N_X3/X14/21_X3/X14/M11_d N_B15_X3/X14/M11_g N_VDD_X3/X14/M11_s
+ N_VDD_X3/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX3/X14/M12 N_X3/X14/13_X3/X14/M12_d N_A15_X3/X14/M12_g N_X3/X14/21_X3/X14/M12_s
+ N_VDD_X3/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX3/X14/M13 N_VDD_X3/X14/M13_d N_X3/X14/13_X3/X14/M13_g N_X3/X14/17_X3/X14/M13_s
+ N_VDD_X3/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X14/X14/M0 N_GND_X3/X14/X14/M0_d N_X3/X14/18_X3/X14/X14/M0_g
+ N_SUM15_X3/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X14/X14/M1 N_X3/X14/X14/10_X3/X14/X14/M1_d N_X3/35_X3/X14/X14/M1_g
+ N_X3/X14/18_X3/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X14/X14/M2 N_GND_X3/X14/X14/M2_d N_X3/29_X3/X14/X14/M2_g
+ N_X3/X14/X14/10_X3/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X14/X14/M3 N_X3/X14/X14/11_X3/X14/X14/M3_d N_X3/X14/16_X3/X14/X14/M3_g
+ N_GND_X3/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X14/X14/M4 N_X3/X14/18_X3/X14/X14/M4_d N_X3/38_X3/X14/X14/M4_g
+ N_X3/X14/X14/11_X3/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X14/X14/M5 N_X3/X14/X14/9_X3/X14/X14/M5_d N_X3/X14/16_X3/X14/X14/M5_g
+ N_VDD_X3/X14/X14/M5_s N_VDD_X3/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X14/X14/M6 N_X3/X14/18_X3/X14/X14/M6_d N_X3/35_X3/X14/X14/M6_g
+ N_X3/X14/X14/9_X3/X14/X14/M6_s N_VDD_X3/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X14/M7 N_X3/X14/X14/9_X3/X14/X14/M7_d N_X3/29_X3/X14/X14/M7_g
+ N_X3/X14/18_X3/X14/X14/M7_s N_VDD_X3/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X14/M8 N_VDD_X3/X14/X14/M8_d N_X3/38_X3/X14/X14/M8_g
+ N_X3/X14/X14/9_X3/X14/X14/M8_s N_VDD_X3/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X14/X14/M9 N_VDD_X3/X14/X14/M9_d N_X3/X14/18_X3/X14/X14/M9_g
+ N_SUM15_X3/X14/X14/M9_s N_VDD_X3/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X14/X15/M0 N_GND_X3/X14/X15/M0_d N_X3/33_X3/X14/X15/M0_g
+ N_X3/34_X3/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X14/X15/M1 N_X3/X14/X15/10_X3/X14/X15/M1_d N_X3/X14/17_X3/X14/X15/M1_g
+ N_X3/33_X3/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX3/X14/X15/M2 N_GND_X3/X14/X15/M2_d N_X3/38_X3/X14/X15/M2_g
+ N_X3/X14/X15/10_X3/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X14/X15/M3 N_X3/X14/X15/11_X3/X14/X15/M3_d N_B15_X3/X14/X15/M3_g
+ N_GND_X3/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X14/X15/M4 N_X3/33_X3/X14/X15/M4_d N_A15_X3/X14/X15/M4_g
+ N_X3/X14/X15/11_X3/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X14/X15/M5 N_X3/X14/X15/9_X3/X14/X15/M5_d N_B15_X3/X14/X15/M5_g
+ N_VDD_X3/X14/X15/M5_s N_VDD_X3/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X14/X15/M6 N_X3/33_X3/X14/X15/M6_d N_X3/X14/17_X3/X14/X15/M6_g
+ N_X3/X14/X15/9_X3/X14/X15/M6_s N_VDD_X3/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X15/M7 N_X3/X14/X15/9_X3/X14/X15/M7_d N_X3/38_X3/X14/X15/M7_g
+ N_X3/33_X3/X14/X15/M7_s N_VDD_X3/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X15/M8 N_VDD_X3/X14/X15/M8_d N_A15_X3/X14/X15/M8_g
+ N_X3/X14/X15/9_X3/X14/X15/M8_s N_VDD_X3/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X14/X15/M9 N_VDD_X3/X14/X15/M9_d N_X3/33_X3/X14/X15/M9_g
+ N_X3/34_X3/X14/X15/M9_s N_VDD_X3/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX3/X14/X16/M0 N_GND_X3/X14/X16/M0_d N_X3/X14/19_X3/X14/X16/M0_g
+ N_X3/35_X3/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX3/X14/X16/M1 N_X3/X14/X16/10_X3/X14/X16/M1_d N_A15N_X3/X14/X16/M1_g
+ N_X3/X14/19_X3/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX3/X14/X16/M2 N_GND_X3/X14/X16/M2_d N_B15_X3/X14/X16/M2_g
+ N_X3/X14/X16/10_X3/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX3/X14/X16/M3 N_X3/X14/X16/11_X3/X14/X16/M3_d N_B15N_X3/X14/X16/M3_g
+ N_GND_X3/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX3/X14/X16/M4 N_X3/X14/19_X3/X14/X16/M4_d N_A15_X3/X14/X16/M4_g
+ N_X3/X14/X16/11_X3/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX3/X14/X16/M5 N_X3/X14/X16/9_X3/X14/X16/M5_d N_B15N_X3/X14/X16/M5_g
+ N_VDD_X3/X14/X16/M5_s N_VDD_X3/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX3/X14/X16/M6 N_X3/X14/19_X3/X14/X16/M6_d N_A15N_X3/X14/X16/M6_g
+ N_X3/X14/X16/9_X3/X14/X16/M6_s N_VDD_X3/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X16/M7 N_X3/X14/X16/9_X3/X14/X16/M7_d N_B15_X3/X14/X16/M7_g
+ N_X3/X14/19_X3/X14/X16/M7_s N_VDD_X3/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX3/X14/X16/M8 N_VDD_X3/X14/X16/M8_d N_A15_X3/X14/X16/M8_g
+ N_X3/X14/X16/9_X3/X14/X16/M8_s N_VDD_X3/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX3/X14/X16/M9 N_VDD_X3/X14/X16/M9_d N_X3/X14/19_X3/X14/X16/M9_g
+ N_X3/35_X3/X14/X16/M9_s N_VDD_X3/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/M0 N_GND_X4/M0_d N_X4/39_X4/M0_g N_X4/40_X4/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/M1 N_X4/41_X4/M1_d N_X4/32_X4/M1_g N_GND_X4/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX4/M2 N_X4/42_X4/M2_d N_X4/31_X4/M2_g N_X4/41_X4/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX4/M3 N_X4/43_X4/M3_d N_X4/30_X4/M3_g N_X4/42_X4/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX4/M4 N_X4/39_X4/M4_d N_X4/35_X4/M4_g N_X4/43_X4/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX4/M5 N_VDD_X4/M5_d N_X4/39_X4/M5_g N_X4/40_X4/M5_s N_VDD_X4/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/M6 N_X4/39_X4/M6_d N_X4/32_X4/M6_g N_VDD_X4/M6_s N_VDD_X4/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX4/M7 N_VDD_X4/M7_d N_X4/31_X4/M7_g N_X4/39_X4/M7_s N_VDD_X4/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX4/M8 N_X4/39_X4/M8_d N_X4/30_X4/M8_g N_VDD_X4/M8_s N_VDD_X4/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX4/M9 N_VDD_X4/M9_d N_X4/35_X4/M9_g N_X4/39_X4/M9_s N_VDD_X4/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX4/X10/M0 N_GND_X4/X10/M0_d N_6_X4/X10/M0_g N_48_X4/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X10/M1 N_X4/X10/10_X4/X10/M1_d N_49_X4/X10/M1_g N_6_X4/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X10/M2 N_GND_X4/X10/M2_d N_X4/40_X4/X10/M2_g N_X4/X10/10_X4/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X10/M3 N_X4/X10/11_X4/X10/M3_d N_X4/39_X4/X10/M3_g N_GND_X4/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X10/M4 N_6_X4/X10/M4_d N_X4/34_X4/X10/M4_g N_X4/X10/11_X4/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X10/M5 N_X4/X10/9_X4/X10/M5_d N_X4/39_X4/X10/M5_g N_VDD_X4/X10/M5_s
+ N_VDD_X4/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX4/X10/M6 N_6_X4/X10/M6_d N_49_X4/X10/M6_g N_X4/X10/9_X4/X10/M6_s
+ N_VDD_X4/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X10/M7 N_X4/X10/9_X4/X10/M7_d N_X4/40_X4/X10/M7_g N_6_X4/X10/M7_s
+ N_VDD_X4/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X10/M8 N_VDD_X4/X10/M8_d N_X4/34_X4/X10/M8_g N_X4/X10/9_X4/X10/M8_s
+ N_VDD_X4/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X10/M9 N_VDD_X4/X10/M9_d N_6_X4/X10/M9_g N_48_X4/X10/M9_s N_VDD_X4/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X11/M0 N_GND_X4/X11/M0_d N_X4/X11/14_X4/X11/M0_g N_X4/X11/16_X4/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X11/M1 N_GND_X4/X11/M1_d N_X4/X11/13_X4/X11/M1_g N_X4/X11/14_X4/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X11/M2 N_X4/X11/20_X4/X11/M2_d N_B10_X4/X11/M2_g N_GND_X4/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X11/M3 N_X4/X11/14_X4/X11/M3_d N_A10_X4/X11/M3_g N_X4/X11/20_X4/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X11/M4 N_GND_X4/X11/M4_d N_X4/X11/13_X4/X11/M4_g N_X4/X11/17_X4/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X11/M5 N_X4/X11/13_X4/X11/M5_d N_B10_X4/X11/M5_g N_GND_X4/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X11/M6 N_GND_X4/X11/M6_d N_A10_X4/X11/M6_g N_X4/X11/13_X4/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X11/M7 N_X4/X11/15_X4/X11/M7_d N_X4/X11/13_X4/X11/M7_g
+ N_X4/X11/14_X4/X11/M7_s N_VDD_X4/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX4/X11/M8 N_VDD_X4/X11/M8_d N_B10_X4/X11/M8_g N_X4/X11/15_X4/X11/M8_s
+ N_VDD_X4/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X11/M9 N_X4/X11/15_X4/X11/M9_d N_A10_X4/X11/M9_g N_VDD_X4/X11/M9_s
+ N_VDD_X4/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X11/M10 N_VDD_X4/X11/M10_d N_X4/X11/14_X4/X11/M10_g N_X4/X11/16_X4/X11/M10_s
+ N_VDD_X4/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X11/M11 N_X4/X11/21_X4/X11/M11_d N_B10_X4/X11/M11_g N_VDD_X4/X11/M11_s
+ N_VDD_X4/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX4/X11/M12 N_X4/X11/13_X4/X11/M12_d N_A10_X4/X11/M12_g N_X4/X11/21_X4/X11/M12_s
+ N_VDD_X4/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X11/M13 N_VDD_X4/X11/M13_d N_X4/X11/13_X4/X11/M13_g N_X4/X11/17_X4/X11/M13_s
+ N_VDD_X4/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X11/X14/M0 N_GND_X4/X11/X14/M0_d N_X4/X11/18_X4/X11/X14/M0_g
+ N_SUM10_X4/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X11/X14/M1 N_X4/X11/X14/10_X4/X11/X14/M1_d N_X4/30_X4/X11/X14/M1_g
+ N_X4/X11/18_X4/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X11/X14/M2 N_GND_X4/X11/X14/M2_d N_X4/27_X4/X11/X14/M2_g
+ N_X4/X11/X14/10_X4/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X11/X14/M3 N_X4/X11/X14/11_X4/X11/X14/M3_d N_X4/X11/16_X4/X11/X14/M3_g
+ N_GND_X4/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X11/X14/M4 N_X4/X11/18_X4/X11/X14/M4_d N_X4/36_X4/X11/X14/M4_g
+ N_X4/X11/X14/11_X4/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X11/X14/M5 N_X4/X11/X14/9_X4/X11/X14/M5_d N_X4/X11/16_X4/X11/X14/M5_g
+ N_VDD_X4/X11/X14/M5_s N_VDD_X4/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X11/X14/M6 N_X4/X11/18_X4/X11/X14/M6_d N_X4/30_X4/X11/X14/M6_g
+ N_X4/X11/X14/9_X4/X11/X14/M6_s N_VDD_X4/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X14/M7 N_X4/X11/X14/9_X4/X11/X14/M7_d N_X4/27_X4/X11/X14/M7_g
+ N_X4/X11/18_X4/X11/X14/M7_s N_VDD_X4/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X14/M8 N_VDD_X4/X11/X14/M8_d N_X4/36_X4/X11/X14/M8_g
+ N_X4/X11/X14/9_X4/X11/X14/M8_s N_VDD_X4/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X11/X14/M9 N_VDD_X4/X11/X14/M9_d N_X4/X11/18_X4/X11/X14/M9_g
+ N_SUM10_X4/X11/X14/M9_s N_VDD_X4/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X11/X15/M0 N_GND_X4/X11/X15/M0_d N_X4/29_X4/X11/X15/M0_g
+ N_X4/38_X4/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X11/X15/M1 N_X4/X11/X15/10_X4/X11/X15/M1_d N_X4/X11/17_X4/X11/X15/M1_g
+ N_X4/29_X4/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX4/X11/X15/M2 N_GND_X4/X11/X15/M2_d N_X4/36_X4/X11/X15/M2_g
+ N_X4/X11/X15/10_X4/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X11/X15/M3 N_X4/X11/X15/11_X4/X11/X15/M3_d N_B10_X4/X11/X15/M3_g
+ N_GND_X4/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X11/X15/M4 N_X4/29_X4/X11/X15/M4_d N_A10_X4/X11/X15/M4_g
+ N_X4/X11/X15/11_X4/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X11/X15/M5 N_X4/X11/X15/9_X4/X11/X15/M5_d N_B10_X4/X11/X15/M5_g
+ N_VDD_X4/X11/X15/M5_s N_VDD_X4/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X11/X15/M6 N_X4/29_X4/X11/X15/M6_d N_X4/X11/17_X4/X11/X15/M6_g
+ N_X4/X11/X15/9_X4/X11/X15/M6_s N_VDD_X4/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X15/M7 N_X4/X11/X15/9_X4/X11/X15/M7_d N_X4/36_X4/X11/X15/M7_g
+ N_X4/29_X4/X11/X15/M7_s N_VDD_X4/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X15/M8 N_VDD_X4/X11/X15/M8_d N_A10_X4/X11/X15/M8_g
+ N_X4/X11/X15/9_X4/X11/X15/M8_s N_VDD_X4/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X11/X15/M9 N_VDD_X4/X11/X15/M9_d N_X4/29_X4/X11/X15/M9_g
+ N_X4/38_X4/X11/X15/M9_s N_VDD_X4/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X11/X16/M0 N_GND_X4/X11/X16/M0_d N_X4/X11/19_X4/X11/X16/M0_g
+ N_X4/30_X4/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X11/X16/M1 N_X4/X11/X16/10_X4/X11/X16/M1_d N_A10N_X4/X11/X16/M1_g
+ N_X4/X11/19_X4/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X11/X16/M2 N_GND_X4/X11/X16/M2_d N_B10_X4/X11/X16/M2_g
+ N_X4/X11/X16/10_X4/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X11/X16/M3 N_X4/X11/X16/11_X4/X11/X16/M3_d N_B10N_X4/X11/X16/M3_g
+ N_GND_X4/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X11/X16/M4 N_X4/X11/19_X4/X11/X16/M4_d N_A10_X4/X11/X16/M4_g
+ N_X4/X11/X16/11_X4/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X11/X16/M5 N_X4/X11/X16/9_X4/X11/X16/M5_d N_B10N_X4/X11/X16/M5_g
+ N_VDD_X4/X11/X16/M5_s N_VDD_X4/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X11/X16/M6 N_X4/X11/19_X4/X11/X16/M6_d N_A10N_X4/X11/X16/M6_g
+ N_X4/X11/X16/9_X4/X11/X16/M6_s N_VDD_X4/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X16/M7 N_X4/X11/X16/9_X4/X11/X16/M7_d N_B10_X4/X11/X16/M7_g
+ N_X4/X11/19_X4/X11/X16/M7_s N_VDD_X4/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X11/X16/M8 N_VDD_X4/X11/X16/M8_d N_A10_X4/X11/X16/M8_g
+ N_X4/X11/X16/9_X4/X11/X16/M8_s N_VDD_X4/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X11/X16/M9 N_VDD_X4/X11/X16/M9_d N_X4/X11/19_X4/X11/X16/M9_g
+ N_X4/30_X4/X11/X16/M9_s N_VDD_X4/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X12/M0 N_GND_X4/X12/M0_d N_X4/X12/14_X4/X12/M0_g N_X4/X12/16_X4/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X12/M1 N_GND_X4/X12/M1_d N_X4/X12/13_X4/X12/M1_g N_X4/X12/14_X4/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X12/M2 N_X4/X12/20_X4/X12/M2_d N_B9_X4/X12/M2_g N_GND_X4/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X12/M3 N_X4/X12/14_X4/X12/M3_d N_A9_X4/X12/M3_g N_X4/X12/20_X4/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X12/M4 N_GND_X4/X12/M4_d N_X4/X12/13_X4/X12/M4_g N_X4/X12/17_X4/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X12/M5 N_X4/X12/13_X4/X12/M5_d N_B9_X4/X12/M5_g N_GND_X4/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X12/M6 N_GND_X4/X12/M6_d N_A9_X4/X12/M6_g N_X4/X12/13_X4/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X12/M7 N_X4/X12/15_X4/X12/M7_d N_X4/X12/13_X4/X12/M7_g
+ N_X4/X12/14_X4/X12/M7_s N_VDD_X4/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX4/X12/M8 N_VDD_X4/X12/M8_d N_B9_X4/X12/M8_g N_X4/X12/15_X4/X12/M8_s
+ N_VDD_X4/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X12/M9 N_X4/X12/15_X4/X12/M9_d N_A9_X4/X12/M9_g N_VDD_X4/X12/M9_s
+ N_VDD_X4/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X12/M10 N_VDD_X4/X12/M10_d N_X4/X12/14_X4/X12/M10_g N_X4/X12/16_X4/X12/M10_s
+ N_VDD_X4/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X12/M11 N_X4/X12/21_X4/X12/M11_d N_B9_X4/X12/M11_g N_VDD_X4/X12/M11_s
+ N_VDD_X4/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX4/X12/M12 N_X4/X12/13_X4/X12/M12_d N_A9_X4/X12/M12_g N_X4/X12/21_X4/X12/M12_s
+ N_VDD_X4/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X12/M13 N_VDD_X4/X12/M13_d N_X4/X12/13_X4/X12/M13_g N_X4/X12/17_X4/X12/M13_s
+ N_VDD_X4/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X12/X14/M0 N_GND_X4/X12/X14/M0_d N_X4/X12/18_X4/X12/X14/M0_g
+ N_SUM9_X4/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X12/X14/M1 N_X4/X12/X14/10_X4/X12/X14/M1_d N_X4/31_X4/X12/X14/M1_g
+ N_X4/X12/18_X4/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X12/X14/M2 N_GND_X4/X12/X14/M2_d N_X4/28_X4/X12/X14/M2_g
+ N_X4/X12/X14/10_X4/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X12/X14/M3 N_X4/X12/X14/11_X4/X12/X14/M3_d N_X4/X12/16_X4/X12/X14/M3_g
+ N_GND_X4/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X12/X14/M4 N_X4/X12/18_X4/X12/X14/M4_d N_X4/37_X4/X12/X14/M4_g
+ N_X4/X12/X14/11_X4/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X12/X14/M5 N_X4/X12/X14/9_X4/X12/X14/M5_d N_X4/X12/16_X4/X12/X14/M5_g
+ N_VDD_X4/X12/X14/M5_s N_VDD_X4/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X12/X14/M6 N_X4/X12/18_X4/X12/X14/M6_d N_X4/31_X4/X12/X14/M6_g
+ N_X4/X12/X14/9_X4/X12/X14/M6_s N_VDD_X4/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X14/M7 N_X4/X12/X14/9_X4/X12/X14/M7_d N_X4/28_X4/X12/X14/M7_g
+ N_X4/X12/18_X4/X12/X14/M7_s N_VDD_X4/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X14/M8 N_VDD_X4/X12/X14/M8_d N_X4/37_X4/X12/X14/M8_g
+ N_X4/X12/X14/9_X4/X12/X14/M8_s N_VDD_X4/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X12/X14/M9 N_VDD_X4/X12/X14/M9_d N_X4/X12/18_X4/X12/X14/M9_g
+ N_SUM9_X4/X12/X14/M9_s N_VDD_X4/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X12/X15/M0 N_GND_X4/X12/X15/M0_d N_X4/27_X4/X12/X15/M0_g
+ N_X4/36_X4/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X12/X15/M1 N_X4/X12/X15/10_X4/X12/X15/M1_d N_X4/X12/17_X4/X12/X15/M1_g
+ N_X4/27_X4/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX4/X12/X15/M2 N_GND_X4/X12/X15/M2_d N_X4/37_X4/X12/X15/M2_g
+ N_X4/X12/X15/10_X4/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X12/X15/M3 N_X4/X12/X15/11_X4/X12/X15/M3_d N_B9_X4/X12/X15/M3_g
+ N_GND_X4/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X12/X15/M4 N_X4/27_X4/X12/X15/M4_d N_A9_X4/X12/X15/M4_g
+ N_X4/X12/X15/11_X4/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X12/X15/M5 N_X4/X12/X15/9_X4/X12/X15/M5_d N_B9_X4/X12/X15/M5_g
+ N_VDD_X4/X12/X15/M5_s N_VDD_X4/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X12/X15/M6 N_X4/27_X4/X12/X15/M6_d N_X4/X12/17_X4/X12/X15/M6_g
+ N_X4/X12/X15/9_X4/X12/X15/M6_s N_VDD_X4/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X15/M7 N_X4/X12/X15/9_X4/X12/X15/M7_d N_X4/37_X4/X12/X15/M7_g
+ N_X4/27_X4/X12/X15/M7_s N_VDD_X4/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X15/M8 N_VDD_X4/X12/X15/M8_d N_A9_X4/X12/X15/M8_g
+ N_X4/X12/X15/9_X4/X12/X15/M8_s N_VDD_X4/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X12/X15/M9 N_VDD_X4/X12/X15/M9_d N_X4/27_X4/X12/X15/M9_g
+ N_X4/36_X4/X12/X15/M9_s N_VDD_X4/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X12/X16/M0 N_GND_X4/X12/X16/M0_d N_X4/X12/19_X4/X12/X16/M0_g
+ N_X4/31_X4/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X12/X16/M1 N_X4/X12/X16/10_X4/X12/X16/M1_d N_A9N_X4/X12/X16/M1_g
+ N_X4/X12/19_X4/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X12/X16/M2 N_GND_X4/X12/X16/M2_d N_B9_X4/X12/X16/M2_g
+ N_X4/X12/X16/10_X4/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X12/X16/M3 N_X4/X12/X16/11_X4/X12/X16/M3_d N_B9N_X4/X12/X16/M3_g
+ N_GND_X4/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X12/X16/M4 N_X4/X12/19_X4/X12/X16/M4_d N_A9_X4/X12/X16/M4_g
+ N_X4/X12/X16/11_X4/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X12/X16/M5 N_X4/X12/X16/9_X4/X12/X16/M5_d N_B9N_X4/X12/X16/M5_g
+ N_VDD_X4/X12/X16/M5_s N_VDD_X4/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X12/X16/M6 N_X4/X12/19_X4/X12/X16/M6_d N_A9N_X4/X12/X16/M6_g
+ N_X4/X12/X16/9_X4/X12/X16/M6_s N_VDD_X4/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X16/M7 N_X4/X12/X16/9_X4/X12/X16/M7_d N_B9_X4/X12/X16/M7_g
+ N_X4/X12/19_X4/X12/X16/M7_s N_VDD_X4/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X12/X16/M8 N_VDD_X4/X12/X16/M8_d N_A9_X4/X12/X16/M8_g
+ N_X4/X12/X16/9_X4/X12/X16/M8_s N_VDD_X4/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X12/X16/M9 N_VDD_X4/X12/X16/M9_d N_X4/X12/19_X4/X12/X16/M9_g
+ N_X4/31_X4/X12/X16/M9_s N_VDD_X4/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X13/M0 N_GND_X4/X13/M0_d N_X4/X13/14_X4/X13/M0_g N_X4/X13/16_X4/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X13/M1 N_GND_X4/X13/M1_d N_X4/X13/13_X4/X13/M1_g N_X4/X13/14_X4/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X13/M2 N_X4/X13/20_X4/X13/M2_d N_B8_X4/X13/M2_g N_GND_X4/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X13/M3 N_X4/X13/14_X4/X13/M3_d N_A8_X4/X13/M3_g N_X4/X13/20_X4/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X13/M4 N_GND_X4/X13/M4_d N_X4/X13/13_X4/X13/M4_g N_X4/X13/17_X4/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X13/M5 N_X4/X13/13_X4/X13/M5_d N_B8_X4/X13/M5_g N_GND_X4/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X13/M6 N_GND_X4/X13/M6_d N_A8_X4/X13/M6_g N_X4/X13/13_X4/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X13/M7 N_X4/X13/15_X4/X13/M7_d N_X4/X13/13_X4/X13/M7_g
+ N_X4/X13/14_X4/X13/M7_s N_VDD_X4/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX4/X13/M8 N_VDD_X4/X13/M8_d N_B8_X4/X13/M8_g N_X4/X13/15_X4/X13/M8_s
+ N_VDD_X4/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X13/M9 N_X4/X13/15_X4/X13/M9_d N_A8_X4/X13/M9_g N_VDD_X4/X13/M9_s
+ N_VDD_X4/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X13/M10 N_VDD_X4/X13/M10_d N_X4/X13/14_X4/X13/M10_g N_X4/X13/16_X4/X13/M10_s
+ N_VDD_X4/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X13/M11 N_X4/X13/21_X4/X13/M11_d N_B8_X4/X13/M11_g N_VDD_X4/X13/M11_s
+ N_VDD_X4/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX4/X13/M12 N_X4/X13/13_X4/X13/M12_d N_A8_X4/X13/M12_g N_X4/X13/21_X4/X13/M12_s
+ N_VDD_X4/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X13/M13 N_VDD_X4/X13/M13_d N_X4/X13/13_X4/X13/M13_g N_X4/X13/17_X4/X13/M13_s
+ N_VDD_X4/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X13/X14/M0 N_GND_X4/X13/X14/M0_d N_X4/X13/18_X4/X13/X14/M0_g
+ N_SUM8_X4/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X13/X14/M1 N_X4/X13/X14/10_X4/X13/X14/M1_d N_X4/32_X4/X13/X14/M1_g
+ N_X4/X13/18_X4/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X13/X14/M2 N_GND_X4/X13/X14/M2_d N_7_X4/X13/X14/M2_g
+ N_X4/X13/X14/10_X4/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X13/X14/M3 N_X4/X13/X14/11_X4/X13/X14/M3_d N_X4/X13/16_X4/X13/X14/M3_g
+ N_GND_X4/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X13/X14/M4 N_X4/X13/18_X4/X13/X14/M4_d N_49_X4/X13/X14/M4_g
+ N_X4/X13/X14/11_X4/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X13/X14/M5 N_X4/X13/X14/9_X4/X13/X14/M5_d N_X4/X13/16_X4/X13/X14/M5_g
+ N_VDD_X4/X13/X14/M5_s N_VDD_X4/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X13/X14/M6 N_X4/X13/18_X4/X13/X14/M6_d N_X4/32_X4/X13/X14/M6_g
+ N_X4/X13/X14/9_X4/X13/X14/M6_s N_VDD_X4/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X14/M7 N_X4/X13/X14/9_X4/X13/X14/M7_d N_7_X4/X13/X14/M7_g
+ N_X4/X13/18_X4/X13/X14/M7_s N_VDD_X4/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X14/M8 N_VDD_X4/X13/X14/M8_d N_49_X4/X13/X14/M8_g
+ N_X4/X13/X14/9_X4/X13/X14/M8_s N_VDD_X4/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X13/X14/M9 N_VDD_X4/X13/X14/M9_d N_X4/X13/18_X4/X13/X14/M9_g
+ N_SUM8_X4/X13/X14/M9_s N_VDD_X4/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X13/X15/M0 N_GND_X4/X13/X15/M0_d N_X4/28_X4/X13/X15/M0_g
+ N_X4/37_X4/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X13/X15/M1 N_X4/X13/X15/10_X4/X13/X15/M1_d N_X4/X13/17_X4/X13/X15/M1_g
+ N_X4/28_X4/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX4/X13/X15/M2 N_GND_X4/X13/X15/M2_d N_49_X4/X13/X15/M2_g
+ N_X4/X13/X15/10_X4/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X13/X15/M3 N_X4/X13/X15/11_X4/X13/X15/M3_d N_B8_X4/X13/X15/M3_g
+ N_GND_X4/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X13/X15/M4 N_X4/28_X4/X13/X15/M4_d N_A8_X4/X13/X15/M4_g
+ N_X4/X13/X15/11_X4/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X13/X15/M5 N_X4/X13/X15/9_X4/X13/X15/M5_d N_B8_X4/X13/X15/M5_g
+ N_VDD_X4/X13/X15/M5_s N_VDD_X4/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X13/X15/M6 N_X4/28_X4/X13/X15/M6_d N_X4/X13/17_X4/X13/X15/M6_g
+ N_X4/X13/X15/9_X4/X13/X15/M6_s N_VDD_X4/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X15/M7 N_X4/X13/X15/9_X4/X13/X15/M7_d N_49_X4/X13/X15/M7_g
+ N_X4/28_X4/X13/X15/M7_s N_VDD_X4/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X15/M8 N_VDD_X4/X13/X15/M8_d N_A8_X4/X13/X15/M8_g
+ N_X4/X13/X15/9_X4/X13/X15/M8_s N_VDD_X4/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X13/X15/M9 N_VDD_X4/X13/X15/M9_d N_X4/28_X4/X13/X15/M9_g
+ N_X4/37_X4/X13/X15/M9_s N_VDD_X4/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X13/X16/M0 N_GND_X4/X13/X16/M0_d N_X4/X13/19_X4/X13/X16/M0_g
+ N_X4/32_X4/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X13/X16/M1 N_X4/X13/X16/10_X4/X13/X16/M1_d N_A8N_X4/X13/X16/M1_g
+ N_X4/X13/19_X4/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X13/X16/M2 N_GND_X4/X13/X16/M2_d N_B8_X4/X13/X16/M2_g
+ N_X4/X13/X16/10_X4/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X13/X16/M3 N_X4/X13/X16/11_X4/X13/X16/M3_d N_B8N_X4/X13/X16/M3_g
+ N_GND_X4/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X13/X16/M4 N_X4/X13/19_X4/X13/X16/M4_d N_A8_X4/X13/X16/M4_g
+ N_X4/X13/X16/11_X4/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X13/X16/M5 N_X4/X13/X16/9_X4/X13/X16/M5_d N_B8N_X4/X13/X16/M5_g
+ N_VDD_X4/X13/X16/M5_s N_VDD_X4/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X13/X16/M6 N_X4/X13/19_X4/X13/X16/M6_d N_A8N_X4/X13/X16/M6_g
+ N_X4/X13/X16/9_X4/X13/X16/M6_s N_VDD_X4/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X16/M7 N_X4/X13/X16/9_X4/X13/X16/M7_d N_B8_X4/X13/X16/M7_g
+ N_X4/X13/19_X4/X13/X16/M7_s N_VDD_X4/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X13/X16/M8 N_VDD_X4/X13/X16/M8_d N_A8_X4/X13/X16/M8_g
+ N_X4/X13/X16/9_X4/X13/X16/M8_s N_VDD_X4/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X13/X16/M9 N_VDD_X4/X13/X16/M9_d N_X4/X13/19_X4/X13/X16/M9_g
+ N_X4/32_X4/X13/X16/M9_s N_VDD_X4/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X14/M0 N_GND_X4/X14/M0_d N_X4/X14/14_X4/X14/M0_g N_X4/X14/16_X4/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X14/M1 N_GND_X4/X14/M1_d N_X4/X14/13_X4/X14/M1_g N_X4/X14/14_X4/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X14/M2 N_X4/X14/20_X4/X14/M2_d N_B11_X4/X14/M2_g N_GND_X4/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX4/X14/M3 N_X4/X14/14_X4/X14/M3_d N_A11_X4/X14/M3_g N_X4/X14/20_X4/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X14/M4 N_GND_X4/X14/M4_d N_X4/X14/13_X4/X14/M4_g N_X4/X14/17_X4/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X14/M5 N_X4/X14/13_X4/X14/M5_d N_B11_X4/X14/M5_g N_GND_X4/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX4/X14/M6 N_GND_X4/X14/M6_d N_A11_X4/X14/M6_g N_X4/X14/13_X4/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX4/X14/M7 N_X4/X14/15_X4/X14/M7_d N_X4/X14/13_X4/X14/M7_g
+ N_X4/X14/14_X4/X14/M7_s N_VDD_X4/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX4/X14/M8 N_VDD_X4/X14/M8_d N_B11_X4/X14/M8_g N_X4/X14/15_X4/X14/M8_s
+ N_VDD_X4/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX4/X14/M9 N_X4/X14/15_X4/X14/M9_d N_A11_X4/X14/M9_g N_VDD_X4/X14/M9_s
+ N_VDD_X4/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X14/M10 N_VDD_X4/X14/M10_d N_X4/X14/14_X4/X14/M10_g N_X4/X14/16_X4/X14/M10_s
+ N_VDD_X4/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X14/M11 N_X4/X14/21_X4/X14/M11_d N_B11_X4/X14/M11_g N_VDD_X4/X14/M11_s
+ N_VDD_X4/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX4/X14/M12 N_X4/X14/13_X4/X14/M12_d N_A11_X4/X14/M12_g N_X4/X14/21_X4/X14/M12_s
+ N_VDD_X4/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX4/X14/M13 N_VDD_X4/X14/M13_d N_X4/X14/13_X4/X14/M13_g N_X4/X14/17_X4/X14/M13_s
+ N_VDD_X4/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X14/X14/M0 N_GND_X4/X14/X14/M0_d N_X4/X14/18_X4/X14/X14/M0_g
+ N_SUM11_X4/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X14/X14/M1 N_X4/X14/X14/10_X4/X14/X14/M1_d N_X4/35_X4/X14/X14/M1_g
+ N_X4/X14/18_X4/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X14/X14/M2 N_GND_X4/X14/X14/M2_d N_X4/29_X4/X14/X14/M2_g
+ N_X4/X14/X14/10_X4/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X14/X14/M3 N_X4/X14/X14/11_X4/X14/X14/M3_d N_X4/X14/16_X4/X14/X14/M3_g
+ N_GND_X4/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X14/X14/M4 N_X4/X14/18_X4/X14/X14/M4_d N_X4/38_X4/X14/X14/M4_g
+ N_X4/X14/X14/11_X4/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X14/X14/M5 N_X4/X14/X14/9_X4/X14/X14/M5_d N_X4/X14/16_X4/X14/X14/M5_g
+ N_VDD_X4/X14/X14/M5_s N_VDD_X4/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X14/X14/M6 N_X4/X14/18_X4/X14/X14/M6_d N_X4/35_X4/X14/X14/M6_g
+ N_X4/X14/X14/9_X4/X14/X14/M6_s N_VDD_X4/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X14/M7 N_X4/X14/X14/9_X4/X14/X14/M7_d N_X4/29_X4/X14/X14/M7_g
+ N_X4/X14/18_X4/X14/X14/M7_s N_VDD_X4/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X14/M8 N_VDD_X4/X14/X14/M8_d N_X4/38_X4/X14/X14/M8_g
+ N_X4/X14/X14/9_X4/X14/X14/M8_s N_VDD_X4/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X14/X14/M9 N_VDD_X4/X14/X14/M9_d N_X4/X14/18_X4/X14/X14/M9_g
+ N_SUM11_X4/X14/X14/M9_s N_VDD_X4/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X14/X15/M0 N_GND_X4/X14/X15/M0_d N_X4/33_X4/X14/X15/M0_g
+ N_X4/34_X4/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X14/X15/M1 N_X4/X14/X15/10_X4/X14/X15/M1_d N_X4/X14/17_X4/X14/X15/M1_g
+ N_X4/33_X4/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX4/X14/X15/M2 N_GND_X4/X14/X15/M2_d N_X4/38_X4/X14/X15/M2_g
+ N_X4/X14/X15/10_X4/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X14/X15/M3 N_X4/X14/X15/11_X4/X14/X15/M3_d N_B11_X4/X14/X15/M3_g
+ N_GND_X4/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X14/X15/M4 N_X4/33_X4/X14/X15/M4_d N_A11_X4/X14/X15/M4_g
+ N_X4/X14/X15/11_X4/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X14/X15/M5 N_X4/X14/X15/9_X4/X14/X15/M5_d N_B11_X4/X14/X15/M5_g
+ N_VDD_X4/X14/X15/M5_s N_VDD_X4/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X14/X15/M6 N_X4/33_X4/X14/X15/M6_d N_X4/X14/17_X4/X14/X15/M6_g
+ N_X4/X14/X15/9_X4/X14/X15/M6_s N_VDD_X4/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X15/M7 N_X4/X14/X15/9_X4/X14/X15/M7_d N_X4/38_X4/X14/X15/M7_g
+ N_X4/33_X4/X14/X15/M7_s N_VDD_X4/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X15/M8 N_VDD_X4/X14/X15/M8_d N_A11_X4/X14/X15/M8_g
+ N_X4/X14/X15/9_X4/X14/X15/M8_s N_VDD_X4/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X14/X15/M9 N_VDD_X4/X14/X15/M9_d N_X4/33_X4/X14/X15/M9_g
+ N_X4/34_X4/X14/X15/M9_s N_VDD_X4/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX4/X14/X16/M0 N_GND_X4/X14/X16/M0_d N_X4/X14/19_X4/X14/X16/M0_g
+ N_X4/35_X4/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX4/X14/X16/M1 N_X4/X14/X16/10_X4/X14/X16/M1_d N_A11N_X4/X14/X16/M1_g
+ N_X4/X14/19_X4/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX4/X14/X16/M2 N_GND_X4/X14/X16/M2_d N_B11_X4/X14/X16/M2_g
+ N_X4/X14/X16/10_X4/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX4/X14/X16/M3 N_X4/X14/X16/11_X4/X14/X16/M3_d N_B11N_X4/X14/X16/M3_g
+ N_GND_X4/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX4/X14/X16/M4 N_X4/X14/19_X4/X14/X16/M4_d N_A11_X4/X14/X16/M4_g
+ N_X4/X14/X16/11_X4/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX4/X14/X16/M5 N_X4/X14/X16/9_X4/X14/X16/M5_d N_B11N_X4/X14/X16/M5_g
+ N_VDD_X4/X14/X16/M5_s N_VDD_X4/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX4/X14/X16/M6 N_X4/X14/19_X4/X14/X16/M6_d N_A11N_X4/X14/X16/M6_g
+ N_X4/X14/X16/9_X4/X14/X16/M6_s N_VDD_X4/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X16/M7 N_X4/X14/X16/9_X4/X14/X16/M7_d N_B11_X4/X14/X16/M7_g
+ N_X4/X14/19_X4/X14/X16/M7_s N_VDD_X4/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX4/X14/X16/M8 N_VDD_X4/X14/X16/M8_d N_A11_X4/X14/X16/M8_g
+ N_X4/X14/X16/9_X4/X14/X16/M8_s N_VDD_X4/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX4/X14/X16/M9 N_VDD_X4/X14/X16/M9_d N_X4/X14/19_X4/X14/X16/M9_g
+ N_X4/35_X4/X14/X16/M9_s N_VDD_X4/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/M0 N_GND_X5/M0_d N_X5/39_X5/M0_g N_X5/40_X5/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/M1 N_X5/41_X5/M1_d N_X5/32_X5/M1_g N_GND_X5/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX5/M2 N_X5/42_X5/M2_d N_X5/31_X5/M2_g N_X5/41_X5/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX5/M3 N_X5/43_X5/M3_d N_X5/30_X5/M3_g N_X5/42_X5/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX5/M4 N_X5/39_X5/M4_d N_X5/35_X5/M4_g N_X5/43_X5/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX5/M5 N_VDD_X5/M5_d N_X5/39_X5/M5_g N_X5/40_X5/M5_s N_VDD_X5/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/M6 N_X5/39_X5/M6_d N_X5/32_X5/M6_g N_VDD_X5/M6_s N_VDD_X5/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX5/M7 N_VDD_X5/M7_d N_X5/31_X5/M7_g N_X5/39_X5/M7_s N_VDD_X5/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX5/M8 N_X5/39_X5/M8_d N_X5/30_X5/M8_g N_VDD_X5/M8_s N_VDD_X5/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX5/M9 N_VDD_X5/M9_d N_X5/35_X5/M9_g N_X5/39_X5/M9_s N_VDD_X5/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX5/X10/M0 N_GND_X5/X10/M0_d N_5_X5/X10/M0_g N_47_X5/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X10/M1 N_X5/X10/10_X5/X10/M1_d N_50_X5/X10/M1_g N_5_X5/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X10/M2 N_GND_X5/X10/M2_d N_X5/40_X5/X10/M2_g N_X5/X10/10_X5/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X10/M3 N_X5/X10/11_X5/X10/M3_d N_X5/39_X5/X10/M3_g N_GND_X5/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X10/M4 N_5_X5/X10/M4_d N_X5/34_X5/X10/M4_g N_X5/X10/11_X5/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X10/M5 N_X5/X10/9_X5/X10/M5_d N_X5/39_X5/X10/M5_g N_VDD_X5/X10/M5_s
+ N_VDD_X5/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX5/X10/M6 N_5_X5/X10/M6_d N_50_X5/X10/M6_g N_X5/X10/9_X5/X10/M6_s
+ N_VDD_X5/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X10/M7 N_X5/X10/9_X5/X10/M7_d N_X5/40_X5/X10/M7_g N_5_X5/X10/M7_s
+ N_VDD_X5/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X10/M8 N_VDD_X5/X10/M8_d N_X5/34_X5/X10/M8_g N_X5/X10/9_X5/X10/M8_s
+ N_VDD_X5/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X10/M9 N_VDD_X5/X10/M9_d N_5_X5/X10/M9_g N_47_X5/X10/M9_s N_VDD_X5/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X11/M0 N_GND_X5/X11/M0_d N_X5/X11/14_X5/X11/M0_g N_X5/X11/16_X5/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X11/M1 N_GND_X5/X11/M1_d N_X5/X11/13_X5/X11/M1_g N_X5/X11/14_X5/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X11/M2 N_X5/X11/20_X5/X11/M2_d N_B18_X5/X11/M2_g N_GND_X5/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X11/M3 N_X5/X11/14_X5/X11/M3_d N_A18_X5/X11/M3_g N_X5/X11/20_X5/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X11/M4 N_GND_X5/X11/M4_d N_X5/X11/13_X5/X11/M4_g N_X5/X11/17_X5/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X11/M5 N_X5/X11/13_X5/X11/M5_d N_B18_X5/X11/M5_g N_GND_X5/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X11/M6 N_GND_X5/X11/M6_d N_A18_X5/X11/M6_g N_X5/X11/13_X5/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X11/M7 N_X5/X11/15_X5/X11/M7_d N_X5/X11/13_X5/X11/M7_g
+ N_X5/X11/14_X5/X11/M7_s N_VDD_X5/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX5/X11/M8 N_VDD_X5/X11/M8_d N_B18_X5/X11/M8_g N_X5/X11/15_X5/X11/M8_s
+ N_VDD_X5/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X11/M9 N_X5/X11/15_X5/X11/M9_d N_A18_X5/X11/M9_g N_VDD_X5/X11/M9_s
+ N_VDD_X5/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X11/M10 N_VDD_X5/X11/M10_d N_X5/X11/14_X5/X11/M10_g N_X5/X11/16_X5/X11/M10_s
+ N_VDD_X5/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X11/M11 N_X5/X11/21_X5/X11/M11_d N_B18_X5/X11/M11_g N_VDD_X5/X11/M11_s
+ N_VDD_X5/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX5/X11/M12 N_X5/X11/13_X5/X11/M12_d N_A18_X5/X11/M12_g N_X5/X11/21_X5/X11/M12_s
+ N_VDD_X5/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X11/M13 N_VDD_X5/X11/M13_d N_X5/X11/13_X5/X11/M13_g N_X5/X11/17_X5/X11/M13_s
+ N_VDD_X5/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X11/X14/M0 N_GND_X5/X11/X14/M0_d N_X5/X11/18_X5/X11/X14/M0_g
+ N_SUM18_X5/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X11/X14/M1 N_X5/X11/X14/10_X5/X11/X14/M1_d N_X5/30_X5/X11/X14/M1_g
+ N_X5/X11/18_X5/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X11/X14/M2 N_GND_X5/X11/X14/M2_d N_X5/27_X5/X11/X14/M2_g
+ N_X5/X11/X14/10_X5/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X11/X14/M3 N_X5/X11/X14/11_X5/X11/X14/M3_d N_X5/X11/16_X5/X11/X14/M3_g
+ N_GND_X5/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X11/X14/M4 N_X5/X11/18_X5/X11/X14/M4_d N_X5/36_X5/X11/X14/M4_g
+ N_X5/X11/X14/11_X5/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X11/X14/M5 N_X5/X11/X14/9_X5/X11/X14/M5_d N_X5/X11/16_X5/X11/X14/M5_g
+ N_VDD_X5/X11/X14/M5_s N_VDD_X5/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X11/X14/M6 N_X5/X11/18_X5/X11/X14/M6_d N_X5/30_X5/X11/X14/M6_g
+ N_X5/X11/X14/9_X5/X11/X14/M6_s N_VDD_X5/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X14/M7 N_X5/X11/X14/9_X5/X11/X14/M7_d N_X5/27_X5/X11/X14/M7_g
+ N_X5/X11/18_X5/X11/X14/M7_s N_VDD_X5/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X14/M8 N_VDD_X5/X11/X14/M8_d N_X5/36_X5/X11/X14/M8_g
+ N_X5/X11/X14/9_X5/X11/X14/M8_s N_VDD_X5/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X11/X14/M9 N_VDD_X5/X11/X14/M9_d N_X5/X11/18_X5/X11/X14/M9_g
+ N_SUM18_X5/X11/X14/M9_s N_VDD_X5/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X11/X15/M0 N_GND_X5/X11/X15/M0_d N_X5/29_X5/X11/X15/M0_g
+ N_X5/38_X5/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X11/X15/M1 N_X5/X11/X15/10_X5/X11/X15/M1_d N_X5/X11/17_X5/X11/X15/M1_g
+ N_X5/29_X5/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX5/X11/X15/M2 N_GND_X5/X11/X15/M2_d N_X5/36_X5/X11/X15/M2_g
+ N_X5/X11/X15/10_X5/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X11/X15/M3 N_X5/X11/X15/11_X5/X11/X15/M3_d N_B18_X5/X11/X15/M3_g
+ N_GND_X5/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X11/X15/M4 N_X5/29_X5/X11/X15/M4_d N_A18_X5/X11/X15/M4_g
+ N_X5/X11/X15/11_X5/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X11/X15/M5 N_X5/X11/X15/9_X5/X11/X15/M5_d N_B18_X5/X11/X15/M5_g
+ N_VDD_X5/X11/X15/M5_s N_VDD_X5/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X11/X15/M6 N_X5/29_X5/X11/X15/M6_d N_X5/X11/17_X5/X11/X15/M6_g
+ N_X5/X11/X15/9_X5/X11/X15/M6_s N_VDD_X5/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X15/M7 N_X5/X11/X15/9_X5/X11/X15/M7_d N_X5/36_X5/X11/X15/M7_g
+ N_X5/29_X5/X11/X15/M7_s N_VDD_X5/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X15/M8 N_VDD_X5/X11/X15/M8_d N_A18_X5/X11/X15/M8_g
+ N_X5/X11/X15/9_X5/X11/X15/M8_s N_VDD_X5/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X11/X15/M9 N_VDD_X5/X11/X15/M9_d N_X5/29_X5/X11/X15/M9_g
+ N_X5/38_X5/X11/X15/M9_s N_VDD_X5/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X11/X16/M0 N_GND_X5/X11/X16/M0_d N_X5/X11/19_X5/X11/X16/M0_g
+ N_X5/30_X5/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X11/X16/M1 N_X5/X11/X16/10_X5/X11/X16/M1_d N_A18N_X5/X11/X16/M1_g
+ N_X5/X11/19_X5/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X11/X16/M2 N_GND_X5/X11/X16/M2_d N_B18_X5/X11/X16/M2_g
+ N_X5/X11/X16/10_X5/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X11/X16/M3 N_X5/X11/X16/11_X5/X11/X16/M3_d N_B18N_X5/X11/X16/M3_g
+ N_GND_X5/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X11/X16/M4 N_X5/X11/19_X5/X11/X16/M4_d N_A18_X5/X11/X16/M4_g
+ N_X5/X11/X16/11_X5/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X11/X16/M5 N_X5/X11/X16/9_X5/X11/X16/M5_d N_B18N_X5/X11/X16/M5_g
+ N_VDD_X5/X11/X16/M5_s N_VDD_X5/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X11/X16/M6 N_X5/X11/19_X5/X11/X16/M6_d N_A18N_X5/X11/X16/M6_g
+ N_X5/X11/X16/9_X5/X11/X16/M6_s N_VDD_X5/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X16/M7 N_X5/X11/X16/9_X5/X11/X16/M7_d N_B18_X5/X11/X16/M7_g
+ N_X5/X11/19_X5/X11/X16/M7_s N_VDD_X5/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X11/X16/M8 N_VDD_X5/X11/X16/M8_d N_A18_X5/X11/X16/M8_g
+ N_X5/X11/X16/9_X5/X11/X16/M8_s N_VDD_X5/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X11/X16/M9 N_VDD_X5/X11/X16/M9_d N_X5/X11/19_X5/X11/X16/M9_g
+ N_X5/30_X5/X11/X16/M9_s N_VDD_X5/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X12/M0 N_GND_X5/X12/M0_d N_X5/X12/14_X5/X12/M0_g N_X5/X12/16_X5/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X12/M1 N_GND_X5/X12/M1_d N_X5/X12/13_X5/X12/M1_g N_X5/X12/14_X5/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X12/M2 N_X5/X12/20_X5/X12/M2_d N_B17_X5/X12/M2_g N_GND_X5/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X12/M3 N_X5/X12/14_X5/X12/M3_d N_A17_X5/X12/M3_g N_X5/X12/20_X5/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X12/M4 N_GND_X5/X12/M4_d N_X5/X12/13_X5/X12/M4_g N_X5/X12/17_X5/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X12/M5 N_X5/X12/13_X5/X12/M5_d N_B17_X5/X12/M5_g N_GND_X5/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X12/M6 N_GND_X5/X12/M6_d N_A17_X5/X12/M6_g N_X5/X12/13_X5/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X12/M7 N_X5/X12/15_X5/X12/M7_d N_X5/X12/13_X5/X12/M7_g
+ N_X5/X12/14_X5/X12/M7_s N_VDD_X5/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX5/X12/M8 N_VDD_X5/X12/M8_d N_B17_X5/X12/M8_g N_X5/X12/15_X5/X12/M8_s
+ N_VDD_X5/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X12/M9 N_X5/X12/15_X5/X12/M9_d N_A17_X5/X12/M9_g N_VDD_X5/X12/M9_s
+ N_VDD_X5/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X12/M10 N_VDD_X5/X12/M10_d N_X5/X12/14_X5/X12/M10_g N_X5/X12/16_X5/X12/M10_s
+ N_VDD_X5/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X12/M11 N_X5/X12/21_X5/X12/M11_d N_B17_X5/X12/M11_g N_VDD_X5/X12/M11_s
+ N_VDD_X5/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX5/X12/M12 N_X5/X12/13_X5/X12/M12_d N_A17_X5/X12/M12_g N_X5/X12/21_X5/X12/M12_s
+ N_VDD_X5/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X12/M13 N_VDD_X5/X12/M13_d N_X5/X12/13_X5/X12/M13_g N_X5/X12/17_X5/X12/M13_s
+ N_VDD_X5/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X12/X14/M0 N_GND_X5/X12/X14/M0_d N_X5/X12/18_X5/X12/X14/M0_g
+ N_SUM17_X5/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X12/X14/M1 N_X5/X12/X14/10_X5/X12/X14/M1_d N_X5/31_X5/X12/X14/M1_g
+ N_X5/X12/18_X5/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X12/X14/M2 N_GND_X5/X12/X14/M2_d N_X5/28_X5/X12/X14/M2_g
+ N_X5/X12/X14/10_X5/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X12/X14/M3 N_X5/X12/X14/11_X5/X12/X14/M3_d N_X5/X12/16_X5/X12/X14/M3_g
+ N_GND_X5/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X12/X14/M4 N_X5/X12/18_X5/X12/X14/M4_d N_X5/37_X5/X12/X14/M4_g
+ N_X5/X12/X14/11_X5/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X12/X14/M5 N_X5/X12/X14/9_X5/X12/X14/M5_d N_X5/X12/16_X5/X12/X14/M5_g
+ N_VDD_X5/X12/X14/M5_s N_VDD_X5/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X12/X14/M6 N_X5/X12/18_X5/X12/X14/M6_d N_X5/31_X5/X12/X14/M6_g
+ N_X5/X12/X14/9_X5/X12/X14/M6_s N_VDD_X5/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X14/M7 N_X5/X12/X14/9_X5/X12/X14/M7_d N_X5/28_X5/X12/X14/M7_g
+ N_X5/X12/18_X5/X12/X14/M7_s N_VDD_X5/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X14/M8 N_VDD_X5/X12/X14/M8_d N_X5/37_X5/X12/X14/M8_g
+ N_X5/X12/X14/9_X5/X12/X14/M8_s N_VDD_X5/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X12/X14/M9 N_VDD_X5/X12/X14/M9_d N_X5/X12/18_X5/X12/X14/M9_g
+ N_SUM17_X5/X12/X14/M9_s N_VDD_X5/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X12/X15/M0 N_GND_X5/X12/X15/M0_d N_X5/27_X5/X12/X15/M0_g
+ N_X5/36_X5/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X12/X15/M1 N_X5/X12/X15/10_X5/X12/X15/M1_d N_X5/X12/17_X5/X12/X15/M1_g
+ N_X5/27_X5/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX5/X12/X15/M2 N_GND_X5/X12/X15/M2_d N_X5/37_X5/X12/X15/M2_g
+ N_X5/X12/X15/10_X5/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X12/X15/M3 N_X5/X12/X15/11_X5/X12/X15/M3_d N_B17_X5/X12/X15/M3_g
+ N_GND_X5/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X12/X15/M4 N_X5/27_X5/X12/X15/M4_d N_A17_X5/X12/X15/M4_g
+ N_X5/X12/X15/11_X5/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X12/X15/M5 N_X5/X12/X15/9_X5/X12/X15/M5_d N_B17_X5/X12/X15/M5_g
+ N_VDD_X5/X12/X15/M5_s N_VDD_X5/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X12/X15/M6 N_X5/27_X5/X12/X15/M6_d N_X5/X12/17_X5/X12/X15/M6_g
+ N_X5/X12/X15/9_X5/X12/X15/M6_s N_VDD_X5/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X15/M7 N_X5/X12/X15/9_X5/X12/X15/M7_d N_X5/37_X5/X12/X15/M7_g
+ N_X5/27_X5/X12/X15/M7_s N_VDD_X5/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X15/M8 N_VDD_X5/X12/X15/M8_d N_A17_X5/X12/X15/M8_g
+ N_X5/X12/X15/9_X5/X12/X15/M8_s N_VDD_X5/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X12/X15/M9 N_VDD_X5/X12/X15/M9_d N_X5/27_X5/X12/X15/M9_g
+ N_X5/36_X5/X12/X15/M9_s N_VDD_X5/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X12/X16/M0 N_GND_X5/X12/X16/M0_d N_X5/X12/19_X5/X12/X16/M0_g
+ N_X5/31_X5/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X12/X16/M1 N_X5/X12/X16/10_X5/X12/X16/M1_d N_A17N_X5/X12/X16/M1_g
+ N_X5/X12/19_X5/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X12/X16/M2 N_GND_X5/X12/X16/M2_d N_B17_X5/X12/X16/M2_g
+ N_X5/X12/X16/10_X5/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X12/X16/M3 N_X5/X12/X16/11_X5/X12/X16/M3_d N_B17N_X5/X12/X16/M3_g
+ N_GND_X5/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X12/X16/M4 N_X5/X12/19_X5/X12/X16/M4_d N_A17_X5/X12/X16/M4_g
+ N_X5/X12/X16/11_X5/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X12/X16/M5 N_X5/X12/X16/9_X5/X12/X16/M5_d N_B17N_X5/X12/X16/M5_g
+ N_VDD_X5/X12/X16/M5_s N_VDD_X5/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X12/X16/M6 N_X5/X12/19_X5/X12/X16/M6_d N_A17N_X5/X12/X16/M6_g
+ N_X5/X12/X16/9_X5/X12/X16/M6_s N_VDD_X5/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X16/M7 N_X5/X12/X16/9_X5/X12/X16/M7_d N_B17_X5/X12/X16/M7_g
+ N_X5/X12/19_X5/X12/X16/M7_s N_VDD_X5/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X12/X16/M8 N_VDD_X5/X12/X16/M8_d N_A17_X5/X12/X16/M8_g
+ N_X5/X12/X16/9_X5/X12/X16/M8_s N_VDD_X5/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X12/X16/M9 N_VDD_X5/X12/X16/M9_d N_X5/X12/19_X5/X12/X16/M9_g
+ N_X5/31_X5/X12/X16/M9_s N_VDD_X5/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X13/M0 N_GND_X5/X13/M0_d N_X5/X13/14_X5/X13/M0_g N_X5/X13/16_X5/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X13/M1 N_GND_X5/X13/M1_d N_X5/X13/13_X5/X13/M1_g N_X5/X13/14_X5/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X13/M2 N_X5/X13/20_X5/X13/M2_d N_B16_X5/X13/M2_g N_GND_X5/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X13/M3 N_X5/X13/14_X5/X13/M3_d N_A16_X5/X13/M3_g N_X5/X13/20_X5/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X13/M4 N_GND_X5/X13/M4_d N_X5/X13/13_X5/X13/M4_g N_X5/X13/17_X5/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X13/M5 N_X5/X13/13_X5/X13/M5_d N_B16_X5/X13/M5_g N_GND_X5/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X13/M6 N_GND_X5/X13/M6_d N_A16_X5/X13/M6_g N_X5/X13/13_X5/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X13/M7 N_X5/X13/15_X5/X13/M7_d N_X5/X13/13_X5/X13/M7_g
+ N_X5/X13/14_X5/X13/M7_s N_VDD_X5/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX5/X13/M8 N_VDD_X5/X13/M8_d N_B16_X5/X13/M8_g N_X5/X13/15_X5/X13/M8_s
+ N_VDD_X5/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X13/M9 N_X5/X13/15_X5/X13/M9_d N_A16_X5/X13/M9_g N_VDD_X5/X13/M9_s
+ N_VDD_X5/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X13/M10 N_VDD_X5/X13/M10_d N_X5/X13/14_X5/X13/M10_g N_X5/X13/16_X5/X13/M10_s
+ N_VDD_X5/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X13/M11 N_X5/X13/21_X5/X13/M11_d N_B16_X5/X13/M11_g N_VDD_X5/X13/M11_s
+ N_VDD_X5/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX5/X13/M12 N_X5/X13/13_X5/X13/M12_d N_A16_X5/X13/M12_g N_X5/X13/21_X5/X13/M12_s
+ N_VDD_X5/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X13/M13 N_VDD_X5/X13/M13_d N_X5/X13/13_X5/X13/M13_g N_X5/X13/17_X5/X13/M13_s
+ N_VDD_X5/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X13/X14/M0 N_GND_X5/X13/X14/M0_d N_X5/X13/18_X5/X13/X14/M0_g
+ N_SUM16_X5/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X13/X14/M1 N_X5/X13/X14/10_X5/X13/X14/M1_d N_X5/32_X5/X13/X14/M1_g
+ N_X5/X13/18_X5/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X13/X14/M2 N_GND_X5/X13/X14/M2_d N_8_X5/X13/X14/M2_g
+ N_X5/X13/X14/10_X5/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X13/X14/M3 N_X5/X13/X14/11_X5/X13/X14/M3_d N_X5/X13/16_X5/X13/X14/M3_g
+ N_GND_X5/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X13/X14/M4 N_X5/X13/18_X5/X13/X14/M4_d N_50_X5/X13/X14/M4_g
+ N_X5/X13/X14/11_X5/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X13/X14/M5 N_X5/X13/X14/9_X5/X13/X14/M5_d N_X5/X13/16_X5/X13/X14/M5_g
+ N_VDD_X5/X13/X14/M5_s N_VDD_X5/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X13/X14/M6 N_X5/X13/18_X5/X13/X14/M6_d N_X5/32_X5/X13/X14/M6_g
+ N_X5/X13/X14/9_X5/X13/X14/M6_s N_VDD_X5/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X14/M7 N_X5/X13/X14/9_X5/X13/X14/M7_d N_8_X5/X13/X14/M7_g
+ N_X5/X13/18_X5/X13/X14/M7_s N_VDD_X5/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X14/M8 N_VDD_X5/X13/X14/M8_d N_50_X5/X13/X14/M8_g
+ N_X5/X13/X14/9_X5/X13/X14/M8_s N_VDD_X5/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X13/X14/M9 N_VDD_X5/X13/X14/M9_d N_X5/X13/18_X5/X13/X14/M9_g
+ N_SUM16_X5/X13/X14/M9_s N_VDD_X5/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X13/X15/M0 N_GND_X5/X13/X15/M0_d N_X5/28_X5/X13/X15/M0_g
+ N_X5/37_X5/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X13/X15/M1 N_X5/X13/X15/10_X5/X13/X15/M1_d N_X5/X13/17_X5/X13/X15/M1_g
+ N_X5/28_X5/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX5/X13/X15/M2 N_GND_X5/X13/X15/M2_d N_50_X5/X13/X15/M2_g
+ N_X5/X13/X15/10_X5/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X13/X15/M3 N_X5/X13/X15/11_X5/X13/X15/M3_d N_B16_X5/X13/X15/M3_g
+ N_GND_X5/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X13/X15/M4 N_X5/28_X5/X13/X15/M4_d N_A16_X5/X13/X15/M4_g
+ N_X5/X13/X15/11_X5/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X13/X15/M5 N_X5/X13/X15/9_X5/X13/X15/M5_d N_B16_X5/X13/X15/M5_g
+ N_VDD_X5/X13/X15/M5_s N_VDD_X5/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X13/X15/M6 N_X5/28_X5/X13/X15/M6_d N_X5/X13/17_X5/X13/X15/M6_g
+ N_X5/X13/X15/9_X5/X13/X15/M6_s N_VDD_X5/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X15/M7 N_X5/X13/X15/9_X5/X13/X15/M7_d N_50_X5/X13/X15/M7_g
+ N_X5/28_X5/X13/X15/M7_s N_VDD_X5/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X15/M8 N_VDD_X5/X13/X15/M8_d N_A16_X5/X13/X15/M8_g
+ N_X5/X13/X15/9_X5/X13/X15/M8_s N_VDD_X5/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X13/X15/M9 N_VDD_X5/X13/X15/M9_d N_X5/28_X5/X13/X15/M9_g
+ N_X5/37_X5/X13/X15/M9_s N_VDD_X5/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X13/X16/M0 N_GND_X5/X13/X16/M0_d N_X5/X13/19_X5/X13/X16/M0_g
+ N_X5/32_X5/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X13/X16/M1 N_X5/X13/X16/10_X5/X13/X16/M1_d N_A16N_X5/X13/X16/M1_g
+ N_X5/X13/19_X5/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X13/X16/M2 N_GND_X5/X13/X16/M2_d N_B16_X5/X13/X16/M2_g
+ N_X5/X13/X16/10_X5/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X13/X16/M3 N_X5/X13/X16/11_X5/X13/X16/M3_d N_B16N_X5/X13/X16/M3_g
+ N_GND_X5/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X13/X16/M4 N_X5/X13/19_X5/X13/X16/M4_d N_A16_X5/X13/X16/M4_g
+ N_X5/X13/X16/11_X5/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X13/X16/M5 N_X5/X13/X16/9_X5/X13/X16/M5_d N_B16N_X5/X13/X16/M5_g
+ N_VDD_X5/X13/X16/M5_s N_VDD_X5/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X13/X16/M6 N_X5/X13/19_X5/X13/X16/M6_d N_A16N_X5/X13/X16/M6_g
+ N_X5/X13/X16/9_X5/X13/X16/M6_s N_VDD_X5/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X16/M7 N_X5/X13/X16/9_X5/X13/X16/M7_d N_B16_X5/X13/X16/M7_g
+ N_X5/X13/19_X5/X13/X16/M7_s N_VDD_X5/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X13/X16/M8 N_VDD_X5/X13/X16/M8_d N_A16_X5/X13/X16/M8_g
+ N_X5/X13/X16/9_X5/X13/X16/M8_s N_VDD_X5/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X13/X16/M9 N_VDD_X5/X13/X16/M9_d N_X5/X13/19_X5/X13/X16/M9_g
+ N_X5/32_X5/X13/X16/M9_s N_VDD_X5/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X14/M0 N_GND_X5/X14/M0_d N_X5/X14/14_X5/X14/M0_g N_X5/X14/16_X5/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X14/M1 N_GND_X5/X14/M1_d N_X5/X14/13_X5/X14/M1_g N_X5/X14/14_X5/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X14/M2 N_X5/X14/20_X5/X14/M2_d N_B19_X5/X14/M2_g N_GND_X5/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX5/X14/M3 N_X5/X14/14_X5/X14/M3_d N_A19_X5/X14/M3_g N_X5/X14/20_X5/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X14/M4 N_GND_X5/X14/M4_d N_X5/X14/13_X5/X14/M4_g N_X5/X14/17_X5/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X14/M5 N_X5/X14/13_X5/X14/M5_d N_B19_X5/X14/M5_g N_GND_X5/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX5/X14/M6 N_GND_X5/X14/M6_d N_A19_X5/X14/M6_g N_X5/X14/13_X5/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX5/X14/M7 N_X5/X14/15_X5/X14/M7_d N_X5/X14/13_X5/X14/M7_g
+ N_X5/X14/14_X5/X14/M7_s N_VDD_X5/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX5/X14/M8 N_VDD_X5/X14/M8_d N_B19_X5/X14/M8_g N_X5/X14/15_X5/X14/M8_s
+ N_VDD_X5/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX5/X14/M9 N_X5/X14/15_X5/X14/M9_d N_A19_X5/X14/M9_g N_VDD_X5/X14/M9_s
+ N_VDD_X5/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X14/M10 N_VDD_X5/X14/M10_d N_X5/X14/14_X5/X14/M10_g N_X5/X14/16_X5/X14/M10_s
+ N_VDD_X5/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X14/M11 N_X5/X14/21_X5/X14/M11_d N_B19_X5/X14/M11_g N_VDD_X5/X14/M11_s
+ N_VDD_X5/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX5/X14/M12 N_X5/X14/13_X5/X14/M12_d N_A19_X5/X14/M12_g N_X5/X14/21_X5/X14/M12_s
+ N_VDD_X5/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX5/X14/M13 N_VDD_X5/X14/M13_d N_X5/X14/13_X5/X14/M13_g N_X5/X14/17_X5/X14/M13_s
+ N_VDD_X5/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X14/X14/M0 N_GND_X5/X14/X14/M0_d N_X5/X14/18_X5/X14/X14/M0_g
+ N_SUM19_X5/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X14/X14/M1 N_X5/X14/X14/10_X5/X14/X14/M1_d N_X5/35_X5/X14/X14/M1_g
+ N_X5/X14/18_X5/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X14/X14/M2 N_GND_X5/X14/X14/M2_d N_X5/29_X5/X14/X14/M2_g
+ N_X5/X14/X14/10_X5/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X14/X14/M3 N_X5/X14/X14/11_X5/X14/X14/M3_d N_X5/X14/16_X5/X14/X14/M3_g
+ N_GND_X5/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X14/X14/M4 N_X5/X14/18_X5/X14/X14/M4_d N_X5/38_X5/X14/X14/M4_g
+ N_X5/X14/X14/11_X5/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X14/X14/M5 N_X5/X14/X14/9_X5/X14/X14/M5_d N_X5/X14/16_X5/X14/X14/M5_g
+ N_VDD_X5/X14/X14/M5_s N_VDD_X5/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X14/X14/M6 N_X5/X14/18_X5/X14/X14/M6_d N_X5/35_X5/X14/X14/M6_g
+ N_X5/X14/X14/9_X5/X14/X14/M6_s N_VDD_X5/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X14/M7 N_X5/X14/X14/9_X5/X14/X14/M7_d N_X5/29_X5/X14/X14/M7_g
+ N_X5/X14/18_X5/X14/X14/M7_s N_VDD_X5/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X14/M8 N_VDD_X5/X14/X14/M8_d N_X5/38_X5/X14/X14/M8_g
+ N_X5/X14/X14/9_X5/X14/X14/M8_s N_VDD_X5/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X14/X14/M9 N_VDD_X5/X14/X14/M9_d N_X5/X14/18_X5/X14/X14/M9_g
+ N_SUM19_X5/X14/X14/M9_s N_VDD_X5/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X14/X15/M0 N_GND_X5/X14/X15/M0_d N_X5/33_X5/X14/X15/M0_g
+ N_X5/34_X5/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X14/X15/M1 N_X5/X14/X15/10_X5/X14/X15/M1_d N_X5/X14/17_X5/X14/X15/M1_g
+ N_X5/33_X5/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX5/X14/X15/M2 N_GND_X5/X14/X15/M2_d N_X5/38_X5/X14/X15/M2_g
+ N_X5/X14/X15/10_X5/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X14/X15/M3 N_X5/X14/X15/11_X5/X14/X15/M3_d N_B19_X5/X14/X15/M3_g
+ N_GND_X5/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X14/X15/M4 N_X5/33_X5/X14/X15/M4_d N_A19_X5/X14/X15/M4_g
+ N_X5/X14/X15/11_X5/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X14/X15/M5 N_X5/X14/X15/9_X5/X14/X15/M5_d N_B19_X5/X14/X15/M5_g
+ N_VDD_X5/X14/X15/M5_s N_VDD_X5/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X14/X15/M6 N_X5/33_X5/X14/X15/M6_d N_X5/X14/17_X5/X14/X15/M6_g
+ N_X5/X14/X15/9_X5/X14/X15/M6_s N_VDD_X5/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X15/M7 N_X5/X14/X15/9_X5/X14/X15/M7_d N_X5/38_X5/X14/X15/M7_g
+ N_X5/33_X5/X14/X15/M7_s N_VDD_X5/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X15/M8 N_VDD_X5/X14/X15/M8_d N_A19_X5/X14/X15/M8_g
+ N_X5/X14/X15/9_X5/X14/X15/M8_s N_VDD_X5/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X14/X15/M9 N_VDD_X5/X14/X15/M9_d N_X5/33_X5/X14/X15/M9_g
+ N_X5/34_X5/X14/X15/M9_s N_VDD_X5/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX5/X14/X16/M0 N_GND_X5/X14/X16/M0_d N_X5/X14/19_X5/X14/X16/M0_g
+ N_X5/35_X5/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX5/X14/X16/M1 N_X5/X14/X16/10_X5/X14/X16/M1_d N_A19N_X5/X14/X16/M1_g
+ N_X5/X14/19_X5/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX5/X14/X16/M2 N_GND_X5/X14/X16/M2_d N_B19_X5/X14/X16/M2_g
+ N_X5/X14/X16/10_X5/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX5/X14/X16/M3 N_X5/X14/X16/11_X5/X14/X16/M3_d N_B19N_X5/X14/X16/M3_g
+ N_GND_X5/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX5/X14/X16/M4 N_X5/X14/19_X5/X14/X16/M4_d N_A19_X5/X14/X16/M4_g
+ N_X5/X14/X16/11_X5/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX5/X14/X16/M5 N_X5/X14/X16/9_X5/X14/X16/M5_d N_B19N_X5/X14/X16/M5_g
+ N_VDD_X5/X14/X16/M5_s N_VDD_X5/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX5/X14/X16/M6 N_X5/X14/19_X5/X14/X16/M6_d N_A19N_X5/X14/X16/M6_g
+ N_X5/X14/X16/9_X5/X14/X16/M6_s N_VDD_X5/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X16/M7 N_X5/X14/X16/9_X5/X14/X16/M7_d N_B19_X5/X14/X16/M7_g
+ N_X5/X14/19_X5/X14/X16/M7_s N_VDD_X5/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX5/X14/X16/M8 N_VDD_X5/X14/X16/M8_d N_A19_X5/X14/X16/M8_g
+ N_X5/X14/X16/9_X5/X14/X16/M8_s N_VDD_X5/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX5/X14/X16/M9 N_VDD_X5/X14/X16/M9_d N_X5/X14/19_X5/X14/X16/M9_g
+ N_X5/35_X5/X14/X16/M9_s N_VDD_X5/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/M0 N_GND_X6/M0_d N_X6/39_X6/M0_g N_X6/40_X6/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/M1 N_X6/41_X6/M1_d N_X6/32_X6/M1_g N_GND_X6/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX6/M2 N_X6/42_X6/M2_d N_X6/31_X6/M2_g N_X6/41_X6/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX6/M3 N_X6/43_X6/M3_d N_X6/30_X6/M3_g N_X6/42_X6/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX6/M4 N_X6/39_X6/M4_d N_X6/35_X6/M4_g N_X6/43_X6/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX6/M5 N_VDD_X6/M5_d N_X6/39_X6/M5_g N_X6/40_X6/M5_s N_VDD_X6/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/M6 N_X6/39_X6/M6_d N_X6/32_X6/M6_g N_VDD_X6/M6_s N_VDD_X6/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX6/M7 N_VDD_X6/M7_d N_X6/31_X6/M7_g N_X6/39_X6/M7_s N_VDD_X6/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX6/M8 N_X6/39_X6/M8_d N_X6/30_X6/M8_g N_VDD_X6/M8_s N_VDD_X6/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX6/M9 N_VDD_X6/M9_d N_X6/35_X6/M9_g N_X6/39_X6/M9_s N_VDD_X6/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX6/X10/M0 N_GND_X6/X10/M0_d N_7_X6/X10/M0_g N_49_X6/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X10/M1 N_X6/X10/10_X6/X10/M1_d N_51_X6/X10/M1_g N_7_X6/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X10/M2 N_GND_X6/X10/M2_d N_X6/40_X6/X10/M2_g N_X6/X10/10_X6/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X10/M3 N_X6/X10/11_X6/X10/M3_d N_X6/39_X6/X10/M3_g N_GND_X6/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X10/M4 N_7_X6/X10/M4_d N_X6/34_X6/X10/M4_g N_X6/X10/11_X6/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X10/M5 N_X6/X10/9_X6/X10/M5_d N_X6/39_X6/X10/M5_g N_VDD_X6/X10/M5_s
+ N_VDD_X6/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX6/X10/M6 N_7_X6/X10/M6_d N_51_X6/X10/M6_g N_X6/X10/9_X6/X10/M6_s
+ N_VDD_X6/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X10/M7 N_X6/X10/9_X6/X10/M7_d N_X6/40_X6/X10/M7_g N_7_X6/X10/M7_s
+ N_VDD_X6/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X10/M8 N_VDD_X6/X10/M8_d N_X6/34_X6/X10/M8_g N_X6/X10/9_X6/X10/M8_s
+ N_VDD_X6/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X10/M9 N_VDD_X6/X10/M9_d N_7_X6/X10/M9_g N_49_X6/X10/M9_s N_VDD_X6/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X11/M0 N_GND_X6/X11/M0_d N_X6/X11/14_X6/X11/M0_g N_X6/X11/16_X6/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X11/M1 N_GND_X6/X11/M1_d N_X6/X11/13_X6/X11/M1_g N_X6/X11/14_X6/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X11/M2 N_X6/X11/20_X6/X11/M2_d N_B6_X6/X11/M2_g N_GND_X6/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X11/M3 N_X6/X11/14_X6/X11/M3_d N_A6_X6/X11/M3_g N_X6/X11/20_X6/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X11/M4 N_GND_X6/X11/M4_d N_X6/X11/13_X6/X11/M4_g N_X6/X11/17_X6/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X11/M5 N_X6/X11/13_X6/X11/M5_d N_B6_X6/X11/M5_g N_GND_X6/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X11/M6 N_GND_X6/X11/M6_d N_A6_X6/X11/M6_g N_X6/X11/13_X6/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X11/M7 N_X6/X11/15_X6/X11/M7_d N_X6/X11/13_X6/X11/M7_g
+ N_X6/X11/14_X6/X11/M7_s N_VDD_X6/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX6/X11/M8 N_VDD_X6/X11/M8_d N_B6_X6/X11/M8_g N_X6/X11/15_X6/X11/M8_s
+ N_VDD_X6/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X11/M9 N_X6/X11/15_X6/X11/M9_d N_A6_X6/X11/M9_g N_VDD_X6/X11/M9_s
+ N_VDD_X6/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X11/M10 N_VDD_X6/X11/M10_d N_X6/X11/14_X6/X11/M10_g N_X6/X11/16_X6/X11/M10_s
+ N_VDD_X6/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X11/M11 N_X6/X11/21_X6/X11/M11_d N_B6_X6/X11/M11_g N_VDD_X6/X11/M11_s
+ N_VDD_X6/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX6/X11/M12 N_X6/X11/13_X6/X11/M12_d N_A6_X6/X11/M12_g N_X6/X11/21_X6/X11/M12_s
+ N_VDD_X6/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X11/M13 N_VDD_X6/X11/M13_d N_X6/X11/13_X6/X11/M13_g N_X6/X11/17_X6/X11/M13_s
+ N_VDD_X6/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X11/X14/M0 N_GND_X6/X11/X14/M0_d N_X6/X11/18_X6/X11/X14/M0_g
+ N_SUM6_X6/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X11/X14/M1 N_X6/X11/X14/10_X6/X11/X14/M1_d N_X6/30_X6/X11/X14/M1_g
+ N_X6/X11/18_X6/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X11/X14/M2 N_GND_X6/X11/X14/M2_d N_X6/27_X6/X11/X14/M2_g
+ N_X6/X11/X14/10_X6/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X11/X14/M3 N_X6/X11/X14/11_X6/X11/X14/M3_d N_X6/X11/16_X6/X11/X14/M3_g
+ N_GND_X6/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X11/X14/M4 N_X6/X11/18_X6/X11/X14/M4_d N_X6/36_X6/X11/X14/M4_g
+ N_X6/X11/X14/11_X6/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X11/X14/M5 N_X6/X11/X14/9_X6/X11/X14/M5_d N_X6/X11/16_X6/X11/X14/M5_g
+ N_VDD_X6/X11/X14/M5_s N_VDD_X6/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X11/X14/M6 N_X6/X11/18_X6/X11/X14/M6_d N_X6/30_X6/X11/X14/M6_g
+ N_X6/X11/X14/9_X6/X11/X14/M6_s N_VDD_X6/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X14/M7 N_X6/X11/X14/9_X6/X11/X14/M7_d N_X6/27_X6/X11/X14/M7_g
+ N_X6/X11/18_X6/X11/X14/M7_s N_VDD_X6/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X14/M8 N_VDD_X6/X11/X14/M8_d N_X6/36_X6/X11/X14/M8_g
+ N_X6/X11/X14/9_X6/X11/X14/M8_s N_VDD_X6/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X11/X14/M9 N_VDD_X6/X11/X14/M9_d N_X6/X11/18_X6/X11/X14/M9_g
+ N_SUM6_X6/X11/X14/M9_s N_VDD_X6/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X11/X15/M0 N_GND_X6/X11/X15/M0_d N_X6/29_X6/X11/X15/M0_g
+ N_X6/38_X6/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X11/X15/M1 N_X6/X11/X15/10_X6/X11/X15/M1_d N_X6/X11/17_X6/X11/X15/M1_g
+ N_X6/29_X6/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX6/X11/X15/M2 N_GND_X6/X11/X15/M2_d N_X6/36_X6/X11/X15/M2_g
+ N_X6/X11/X15/10_X6/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X11/X15/M3 N_X6/X11/X15/11_X6/X11/X15/M3_d N_B6_X6/X11/X15/M3_g
+ N_GND_X6/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X11/X15/M4 N_X6/29_X6/X11/X15/M4_d N_A6_X6/X11/X15/M4_g
+ N_X6/X11/X15/11_X6/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X11/X15/M5 N_X6/X11/X15/9_X6/X11/X15/M5_d N_B6_X6/X11/X15/M5_g
+ N_VDD_X6/X11/X15/M5_s N_VDD_X6/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X11/X15/M6 N_X6/29_X6/X11/X15/M6_d N_X6/X11/17_X6/X11/X15/M6_g
+ N_X6/X11/X15/9_X6/X11/X15/M6_s N_VDD_X6/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X15/M7 N_X6/X11/X15/9_X6/X11/X15/M7_d N_X6/36_X6/X11/X15/M7_g
+ N_X6/29_X6/X11/X15/M7_s N_VDD_X6/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X15/M8 N_VDD_X6/X11/X15/M8_d N_A6_X6/X11/X15/M8_g
+ N_X6/X11/X15/9_X6/X11/X15/M8_s N_VDD_X6/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X11/X15/M9 N_VDD_X6/X11/X15/M9_d N_X6/29_X6/X11/X15/M9_g
+ N_X6/38_X6/X11/X15/M9_s N_VDD_X6/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X11/X16/M0 N_GND_X6/X11/X16/M0_d N_X6/X11/19_X6/X11/X16/M0_g
+ N_X6/30_X6/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X11/X16/M1 N_X6/X11/X16/10_X6/X11/X16/M1_d N_A6N_X6/X11/X16/M1_g
+ N_X6/X11/19_X6/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X11/X16/M2 N_GND_X6/X11/X16/M2_d N_B6_X6/X11/X16/M2_g
+ N_X6/X11/X16/10_X6/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X11/X16/M3 N_X6/X11/X16/11_X6/X11/X16/M3_d N_B6N_X6/X11/X16/M3_g
+ N_GND_X6/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X11/X16/M4 N_X6/X11/19_X6/X11/X16/M4_d N_A6_X6/X11/X16/M4_g
+ N_X6/X11/X16/11_X6/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X11/X16/M5 N_X6/X11/X16/9_X6/X11/X16/M5_d N_B6N_X6/X11/X16/M5_g
+ N_VDD_X6/X11/X16/M5_s N_VDD_X6/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X11/X16/M6 N_X6/X11/19_X6/X11/X16/M6_d N_A6N_X6/X11/X16/M6_g
+ N_X6/X11/X16/9_X6/X11/X16/M6_s N_VDD_X6/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X16/M7 N_X6/X11/X16/9_X6/X11/X16/M7_d N_B6_X6/X11/X16/M7_g
+ N_X6/X11/19_X6/X11/X16/M7_s N_VDD_X6/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X11/X16/M8 N_VDD_X6/X11/X16/M8_d N_A6_X6/X11/X16/M8_g
+ N_X6/X11/X16/9_X6/X11/X16/M8_s N_VDD_X6/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X11/X16/M9 N_VDD_X6/X11/X16/M9_d N_X6/X11/19_X6/X11/X16/M9_g
+ N_X6/30_X6/X11/X16/M9_s N_VDD_X6/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X12/M0 N_GND_X6/X12/M0_d N_X6/X12/14_X6/X12/M0_g N_X6/X12/16_X6/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X12/M1 N_GND_X6/X12/M1_d N_X6/X12/13_X6/X12/M1_g N_X6/X12/14_X6/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X12/M2 N_X6/X12/20_X6/X12/M2_d N_B5_X6/X12/M2_g N_GND_X6/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X12/M3 N_X6/X12/14_X6/X12/M3_d N_A5_X6/X12/M3_g N_X6/X12/20_X6/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X12/M4 N_GND_X6/X12/M4_d N_X6/X12/13_X6/X12/M4_g N_X6/X12/17_X6/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X12/M5 N_X6/X12/13_X6/X12/M5_d N_B5_X6/X12/M5_g N_GND_X6/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X12/M6 N_GND_X6/X12/M6_d N_A5_X6/X12/M6_g N_X6/X12/13_X6/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X12/M7 N_X6/X12/15_X6/X12/M7_d N_X6/X12/13_X6/X12/M7_g
+ N_X6/X12/14_X6/X12/M7_s N_VDD_X6/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX6/X12/M8 N_VDD_X6/X12/M8_d N_B5_X6/X12/M8_g N_X6/X12/15_X6/X12/M8_s
+ N_VDD_X6/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X12/M9 N_X6/X12/15_X6/X12/M9_d N_A5_X6/X12/M9_g N_VDD_X6/X12/M9_s
+ N_VDD_X6/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X12/M10 N_VDD_X6/X12/M10_d N_X6/X12/14_X6/X12/M10_g N_X6/X12/16_X6/X12/M10_s
+ N_VDD_X6/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X12/M11 N_X6/X12/21_X6/X12/M11_d N_B5_X6/X12/M11_g N_VDD_X6/X12/M11_s
+ N_VDD_X6/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX6/X12/M12 N_X6/X12/13_X6/X12/M12_d N_A5_X6/X12/M12_g N_X6/X12/21_X6/X12/M12_s
+ N_VDD_X6/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X12/M13 N_VDD_X6/X12/M13_d N_X6/X12/13_X6/X12/M13_g N_X6/X12/17_X6/X12/M13_s
+ N_VDD_X6/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X12/X14/M0 N_GND_X6/X12/X14/M0_d N_X6/X12/18_X6/X12/X14/M0_g
+ N_SUM5_X6/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X12/X14/M1 N_X6/X12/X14/10_X6/X12/X14/M1_d N_X6/31_X6/X12/X14/M1_g
+ N_X6/X12/18_X6/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X12/X14/M2 N_GND_X6/X12/X14/M2_d N_X6/28_X6/X12/X14/M2_g
+ N_X6/X12/X14/10_X6/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X12/X14/M3 N_X6/X12/X14/11_X6/X12/X14/M3_d N_X6/X12/16_X6/X12/X14/M3_g
+ N_GND_X6/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X12/X14/M4 N_X6/X12/18_X6/X12/X14/M4_d N_X6/37_X6/X12/X14/M4_g
+ N_X6/X12/X14/11_X6/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X12/X14/M5 N_X6/X12/X14/9_X6/X12/X14/M5_d N_X6/X12/16_X6/X12/X14/M5_g
+ N_VDD_X6/X12/X14/M5_s N_VDD_X6/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X12/X14/M6 N_X6/X12/18_X6/X12/X14/M6_d N_X6/31_X6/X12/X14/M6_g
+ N_X6/X12/X14/9_X6/X12/X14/M6_s N_VDD_X6/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X14/M7 N_X6/X12/X14/9_X6/X12/X14/M7_d N_X6/28_X6/X12/X14/M7_g
+ N_X6/X12/18_X6/X12/X14/M7_s N_VDD_X6/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X14/M8 N_VDD_X6/X12/X14/M8_d N_X6/37_X6/X12/X14/M8_g
+ N_X6/X12/X14/9_X6/X12/X14/M8_s N_VDD_X6/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X12/X14/M9 N_VDD_X6/X12/X14/M9_d N_X6/X12/18_X6/X12/X14/M9_g
+ N_SUM5_X6/X12/X14/M9_s N_VDD_X6/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X12/X15/M0 N_GND_X6/X12/X15/M0_d N_X6/27_X6/X12/X15/M0_g
+ N_X6/36_X6/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X12/X15/M1 N_X6/X12/X15/10_X6/X12/X15/M1_d N_X6/X12/17_X6/X12/X15/M1_g
+ N_X6/27_X6/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX6/X12/X15/M2 N_GND_X6/X12/X15/M2_d N_X6/37_X6/X12/X15/M2_g
+ N_X6/X12/X15/10_X6/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X12/X15/M3 N_X6/X12/X15/11_X6/X12/X15/M3_d N_B5_X6/X12/X15/M3_g
+ N_GND_X6/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X12/X15/M4 N_X6/27_X6/X12/X15/M4_d N_A5_X6/X12/X15/M4_g
+ N_X6/X12/X15/11_X6/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X12/X15/M5 N_X6/X12/X15/9_X6/X12/X15/M5_d N_B5_X6/X12/X15/M5_g
+ N_VDD_X6/X12/X15/M5_s N_VDD_X6/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X12/X15/M6 N_X6/27_X6/X12/X15/M6_d N_X6/X12/17_X6/X12/X15/M6_g
+ N_X6/X12/X15/9_X6/X12/X15/M6_s N_VDD_X6/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X15/M7 N_X6/X12/X15/9_X6/X12/X15/M7_d N_X6/37_X6/X12/X15/M7_g
+ N_X6/27_X6/X12/X15/M7_s N_VDD_X6/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X15/M8 N_VDD_X6/X12/X15/M8_d N_A5_X6/X12/X15/M8_g
+ N_X6/X12/X15/9_X6/X12/X15/M8_s N_VDD_X6/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X12/X15/M9 N_VDD_X6/X12/X15/M9_d N_X6/27_X6/X12/X15/M9_g
+ N_X6/36_X6/X12/X15/M9_s N_VDD_X6/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X12/X16/M0 N_GND_X6/X12/X16/M0_d N_X6/X12/19_X6/X12/X16/M0_g
+ N_X6/31_X6/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X12/X16/M1 N_X6/X12/X16/10_X6/X12/X16/M1_d N_A5N_X6/X12/X16/M1_g
+ N_X6/X12/19_X6/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X12/X16/M2 N_GND_X6/X12/X16/M2_d N_B5_X6/X12/X16/M2_g
+ N_X6/X12/X16/10_X6/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X12/X16/M3 N_X6/X12/X16/11_X6/X12/X16/M3_d N_B5N_X6/X12/X16/M3_g
+ N_GND_X6/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X12/X16/M4 N_X6/X12/19_X6/X12/X16/M4_d N_A5_X6/X12/X16/M4_g
+ N_X6/X12/X16/11_X6/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X12/X16/M5 N_X6/X12/X16/9_X6/X12/X16/M5_d N_B5N_X6/X12/X16/M5_g
+ N_VDD_X6/X12/X16/M5_s N_VDD_X6/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X12/X16/M6 N_X6/X12/19_X6/X12/X16/M6_d N_A5N_X6/X12/X16/M6_g
+ N_X6/X12/X16/9_X6/X12/X16/M6_s N_VDD_X6/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X16/M7 N_X6/X12/X16/9_X6/X12/X16/M7_d N_B5_X6/X12/X16/M7_g
+ N_X6/X12/19_X6/X12/X16/M7_s N_VDD_X6/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X12/X16/M8 N_VDD_X6/X12/X16/M8_d N_A5_X6/X12/X16/M8_g
+ N_X6/X12/X16/9_X6/X12/X16/M8_s N_VDD_X6/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X12/X16/M9 N_VDD_X6/X12/X16/M9_d N_X6/X12/19_X6/X12/X16/M9_g
+ N_X6/31_X6/X12/X16/M9_s N_VDD_X6/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X13/M0 N_GND_X6/X13/M0_d N_X6/X13/14_X6/X13/M0_g N_X6/X13/16_X6/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X13/M1 N_GND_X6/X13/M1_d N_X6/X13/13_X6/X13/M1_g N_X6/X13/14_X6/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X13/M2 N_X6/X13/20_X6/X13/M2_d N_B4_X6/X13/M2_g N_GND_X6/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X13/M3 N_X6/X13/14_X6/X13/M3_d N_A4_X6/X13/M3_g N_X6/X13/20_X6/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X13/M4 N_GND_X6/X13/M4_d N_X6/X13/13_X6/X13/M4_g N_X6/X13/17_X6/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X13/M5 N_X6/X13/13_X6/X13/M5_d N_B4_X6/X13/M5_g N_GND_X6/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X13/M6 N_GND_X6/X13/M6_d N_A4_X6/X13/M6_g N_X6/X13/13_X6/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X13/M7 N_X6/X13/15_X6/X13/M7_d N_X6/X13/13_X6/X13/M7_g
+ N_X6/X13/14_X6/X13/M7_s N_VDD_X6/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX6/X13/M8 N_VDD_X6/X13/M8_d N_B4_X6/X13/M8_g N_X6/X13/15_X6/X13/M8_s
+ N_VDD_X6/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X13/M9 N_X6/X13/15_X6/X13/M9_d N_A4_X6/X13/M9_g N_VDD_X6/X13/M9_s
+ N_VDD_X6/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X13/M10 N_VDD_X6/X13/M10_d N_X6/X13/14_X6/X13/M10_g N_X6/X13/16_X6/X13/M10_s
+ N_VDD_X6/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X13/M11 N_X6/X13/21_X6/X13/M11_d N_B4_X6/X13/M11_g N_VDD_X6/X13/M11_s
+ N_VDD_X6/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX6/X13/M12 N_X6/X13/13_X6/X13/M12_d N_A4_X6/X13/M12_g N_X6/X13/21_X6/X13/M12_s
+ N_VDD_X6/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X13/M13 N_VDD_X6/X13/M13_d N_X6/X13/13_X6/X13/M13_g N_X6/X13/17_X6/X13/M13_s
+ N_VDD_X6/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X13/X14/M0 N_GND_X6/X13/X14/M0_d N_X6/X13/18_X6/X13/X14/M0_g
+ N_SUM4_X6/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X13/X14/M1 N_X6/X13/X14/10_X6/X13/X14/M1_d N_X6/32_X6/X13/X14/M1_g
+ N_X6/X13/18_X6/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X13/X14/M2 N_GND_X6/X13/X14/M2_d N_9_X6/X13/X14/M2_g
+ N_X6/X13/X14/10_X6/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X13/X14/M3 N_X6/X13/X14/11_X6/X13/X14/M3_d N_X6/X13/16_X6/X13/X14/M3_g
+ N_GND_X6/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X13/X14/M4 N_X6/X13/18_X6/X13/X14/M4_d N_51_X6/X13/X14/M4_g
+ N_X6/X13/X14/11_X6/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X13/X14/M5 N_X6/X13/X14/9_X6/X13/X14/M5_d N_X6/X13/16_X6/X13/X14/M5_g
+ N_VDD_X6/X13/X14/M5_s N_VDD_X6/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X13/X14/M6 N_X6/X13/18_X6/X13/X14/M6_d N_X6/32_X6/X13/X14/M6_g
+ N_X6/X13/X14/9_X6/X13/X14/M6_s N_VDD_X6/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X14/M7 N_X6/X13/X14/9_X6/X13/X14/M7_d N_9_X6/X13/X14/M7_g
+ N_X6/X13/18_X6/X13/X14/M7_s N_VDD_X6/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X14/M8 N_VDD_X6/X13/X14/M8_d N_51_X6/X13/X14/M8_g
+ N_X6/X13/X14/9_X6/X13/X14/M8_s N_VDD_X6/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X13/X14/M9 N_VDD_X6/X13/X14/M9_d N_X6/X13/18_X6/X13/X14/M9_g
+ N_SUM4_X6/X13/X14/M9_s N_VDD_X6/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X13/X15/M0 N_GND_X6/X13/X15/M0_d N_X6/28_X6/X13/X15/M0_g
+ N_X6/37_X6/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X13/X15/M1 N_X6/X13/X15/10_X6/X13/X15/M1_d N_X6/X13/17_X6/X13/X15/M1_g
+ N_X6/28_X6/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX6/X13/X15/M2 N_GND_X6/X13/X15/M2_d N_51_X6/X13/X15/M2_g
+ N_X6/X13/X15/10_X6/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X13/X15/M3 N_X6/X13/X15/11_X6/X13/X15/M3_d N_B4_X6/X13/X15/M3_g
+ N_GND_X6/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X13/X15/M4 N_X6/28_X6/X13/X15/M4_d N_A4_X6/X13/X15/M4_g
+ N_X6/X13/X15/11_X6/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X13/X15/M5 N_X6/X13/X15/9_X6/X13/X15/M5_d N_B4_X6/X13/X15/M5_g
+ N_VDD_X6/X13/X15/M5_s N_VDD_X6/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X13/X15/M6 N_X6/28_X6/X13/X15/M6_d N_X6/X13/17_X6/X13/X15/M6_g
+ N_X6/X13/X15/9_X6/X13/X15/M6_s N_VDD_X6/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X15/M7 N_X6/X13/X15/9_X6/X13/X15/M7_d N_51_X6/X13/X15/M7_g
+ N_X6/28_X6/X13/X15/M7_s N_VDD_X6/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X15/M8 N_VDD_X6/X13/X15/M8_d N_A4_X6/X13/X15/M8_g
+ N_X6/X13/X15/9_X6/X13/X15/M8_s N_VDD_X6/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X13/X15/M9 N_VDD_X6/X13/X15/M9_d N_X6/28_X6/X13/X15/M9_g
+ N_X6/37_X6/X13/X15/M9_s N_VDD_X6/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X13/X16/M0 N_GND_X6/X13/X16/M0_d N_X6/X13/19_X6/X13/X16/M0_g
+ N_X6/32_X6/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X13/X16/M1 N_X6/X13/X16/10_X6/X13/X16/M1_d N_A4N_X6/X13/X16/M1_g
+ N_X6/X13/19_X6/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X13/X16/M2 N_GND_X6/X13/X16/M2_d N_B4_X6/X13/X16/M2_g
+ N_X6/X13/X16/10_X6/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X13/X16/M3 N_X6/X13/X16/11_X6/X13/X16/M3_d N_B4N_X6/X13/X16/M3_g
+ N_GND_X6/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X13/X16/M4 N_X6/X13/19_X6/X13/X16/M4_d N_A4_X6/X13/X16/M4_g
+ N_X6/X13/X16/11_X6/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X13/X16/M5 N_X6/X13/X16/9_X6/X13/X16/M5_d N_B4N_X6/X13/X16/M5_g
+ N_VDD_X6/X13/X16/M5_s N_VDD_X6/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X13/X16/M6 N_X6/X13/19_X6/X13/X16/M6_d N_A4N_X6/X13/X16/M6_g
+ N_X6/X13/X16/9_X6/X13/X16/M6_s N_VDD_X6/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X16/M7 N_X6/X13/X16/9_X6/X13/X16/M7_d N_B4_X6/X13/X16/M7_g
+ N_X6/X13/19_X6/X13/X16/M7_s N_VDD_X6/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X13/X16/M8 N_VDD_X6/X13/X16/M8_d N_A4_X6/X13/X16/M8_g
+ N_X6/X13/X16/9_X6/X13/X16/M8_s N_VDD_X6/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X13/X16/M9 N_VDD_X6/X13/X16/M9_d N_X6/X13/19_X6/X13/X16/M9_g
+ N_X6/32_X6/X13/X16/M9_s N_VDD_X6/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X14/M0 N_GND_X6/X14/M0_d N_X6/X14/14_X6/X14/M0_g N_X6/X14/16_X6/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X14/M1 N_GND_X6/X14/M1_d N_X6/X14/13_X6/X14/M1_g N_X6/X14/14_X6/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X14/M2 N_X6/X14/20_X6/X14/M2_d N_B7_X6/X14/M2_g N_GND_X6/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX6/X14/M3 N_X6/X14/14_X6/X14/M3_d N_A7_X6/X14/M3_g N_X6/X14/20_X6/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X14/M4 N_GND_X6/X14/M4_d N_X6/X14/13_X6/X14/M4_g N_X6/X14/17_X6/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X14/M5 N_X6/X14/13_X6/X14/M5_d N_B7_X6/X14/M5_g N_GND_X6/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX6/X14/M6 N_GND_X6/X14/M6_d N_A7_X6/X14/M6_g N_X6/X14/13_X6/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX6/X14/M7 N_X6/X14/15_X6/X14/M7_d N_X6/X14/13_X6/X14/M7_g
+ N_X6/X14/14_X6/X14/M7_s N_VDD_X6/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX6/X14/M8 N_VDD_X6/X14/M8_d N_B7_X6/X14/M8_g N_X6/X14/15_X6/X14/M8_s
+ N_VDD_X6/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX6/X14/M9 N_X6/X14/15_X6/X14/M9_d N_A7_X6/X14/M9_g N_VDD_X6/X14/M9_s
+ N_VDD_X6/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X14/M10 N_VDD_X6/X14/M10_d N_X6/X14/14_X6/X14/M10_g N_X6/X14/16_X6/X14/M10_s
+ N_VDD_X6/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X14/M11 N_X6/X14/21_X6/X14/M11_d N_B7_X6/X14/M11_g N_VDD_X6/X14/M11_s
+ N_VDD_X6/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX6/X14/M12 N_X6/X14/13_X6/X14/M12_d N_A7_X6/X14/M12_g N_X6/X14/21_X6/X14/M12_s
+ N_VDD_X6/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX6/X14/M13 N_VDD_X6/X14/M13_d N_X6/X14/13_X6/X14/M13_g N_X6/X14/17_X6/X14/M13_s
+ N_VDD_X6/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X14/X14/M0 N_GND_X6/X14/X14/M0_d N_X6/X14/18_X6/X14/X14/M0_g
+ N_SUM7_X6/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X14/X14/M1 N_X6/X14/X14/10_X6/X14/X14/M1_d N_X6/35_X6/X14/X14/M1_g
+ N_X6/X14/18_X6/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X14/X14/M2 N_GND_X6/X14/X14/M2_d N_X6/29_X6/X14/X14/M2_g
+ N_X6/X14/X14/10_X6/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X14/X14/M3 N_X6/X14/X14/11_X6/X14/X14/M3_d N_X6/X14/16_X6/X14/X14/M3_g
+ N_GND_X6/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X14/X14/M4 N_X6/X14/18_X6/X14/X14/M4_d N_X6/38_X6/X14/X14/M4_g
+ N_X6/X14/X14/11_X6/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X14/X14/M5 N_X6/X14/X14/9_X6/X14/X14/M5_d N_X6/X14/16_X6/X14/X14/M5_g
+ N_VDD_X6/X14/X14/M5_s N_VDD_X6/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X14/X14/M6 N_X6/X14/18_X6/X14/X14/M6_d N_X6/35_X6/X14/X14/M6_g
+ N_X6/X14/X14/9_X6/X14/X14/M6_s N_VDD_X6/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X14/M7 N_X6/X14/X14/9_X6/X14/X14/M7_d N_X6/29_X6/X14/X14/M7_g
+ N_X6/X14/18_X6/X14/X14/M7_s N_VDD_X6/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X14/M8 N_VDD_X6/X14/X14/M8_d N_X6/38_X6/X14/X14/M8_g
+ N_X6/X14/X14/9_X6/X14/X14/M8_s N_VDD_X6/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X14/X14/M9 N_VDD_X6/X14/X14/M9_d N_X6/X14/18_X6/X14/X14/M9_g
+ N_SUM7_X6/X14/X14/M9_s N_VDD_X6/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X14/X15/M0 N_GND_X6/X14/X15/M0_d N_X6/33_X6/X14/X15/M0_g
+ N_X6/34_X6/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X14/X15/M1 N_X6/X14/X15/10_X6/X14/X15/M1_d N_X6/X14/17_X6/X14/X15/M1_g
+ N_X6/33_X6/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX6/X14/X15/M2 N_GND_X6/X14/X15/M2_d N_X6/38_X6/X14/X15/M2_g
+ N_X6/X14/X15/10_X6/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X14/X15/M3 N_X6/X14/X15/11_X6/X14/X15/M3_d N_B7_X6/X14/X15/M3_g
+ N_GND_X6/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X14/X15/M4 N_X6/33_X6/X14/X15/M4_d N_A7_X6/X14/X15/M4_g
+ N_X6/X14/X15/11_X6/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X14/X15/M5 N_X6/X14/X15/9_X6/X14/X15/M5_d N_B7_X6/X14/X15/M5_g
+ N_VDD_X6/X14/X15/M5_s N_VDD_X6/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X14/X15/M6 N_X6/33_X6/X14/X15/M6_d N_X6/X14/17_X6/X14/X15/M6_g
+ N_X6/X14/X15/9_X6/X14/X15/M6_s N_VDD_X6/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X15/M7 N_X6/X14/X15/9_X6/X14/X15/M7_d N_X6/38_X6/X14/X15/M7_g
+ N_X6/33_X6/X14/X15/M7_s N_VDD_X6/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X15/M8 N_VDD_X6/X14/X15/M8_d N_A7_X6/X14/X15/M8_g
+ N_X6/X14/X15/9_X6/X14/X15/M8_s N_VDD_X6/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X14/X15/M9 N_VDD_X6/X14/X15/M9_d N_X6/33_X6/X14/X15/M9_g
+ N_X6/34_X6/X14/X15/M9_s N_VDD_X6/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX6/X14/X16/M0 N_GND_X6/X14/X16/M0_d N_X6/X14/19_X6/X14/X16/M0_g
+ N_X6/35_X6/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX6/X14/X16/M1 N_X6/X14/X16/10_X6/X14/X16/M1_d N_A7N_X6/X14/X16/M1_g
+ N_X6/X14/19_X6/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX6/X14/X16/M2 N_GND_X6/X14/X16/M2_d N_B7_X6/X14/X16/M2_g
+ N_X6/X14/X16/10_X6/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX6/X14/X16/M3 N_X6/X14/X16/11_X6/X14/X16/M3_d N_B7N_X6/X14/X16/M3_g
+ N_GND_X6/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX6/X14/X16/M4 N_X6/X14/19_X6/X14/X16/M4_d N_A7_X6/X14/X16/M4_g
+ N_X6/X14/X16/11_X6/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX6/X14/X16/M5 N_X6/X14/X16/9_X6/X14/X16/M5_d N_B7N_X6/X14/X16/M5_g
+ N_VDD_X6/X14/X16/M5_s N_VDD_X6/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX6/X14/X16/M6 N_X6/X14/19_X6/X14/X16/M6_d N_A7N_X6/X14/X16/M6_g
+ N_X6/X14/X16/9_X6/X14/X16/M6_s N_VDD_X6/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X16/M7 N_X6/X14/X16/9_X6/X14/X16/M7_d N_B7_X6/X14/X16/M7_g
+ N_X6/X14/19_X6/X14/X16/M7_s N_VDD_X6/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX6/X14/X16/M8 N_VDD_X6/X14/X16/M8_d N_A7_X6/X14/X16/M8_g
+ N_X6/X14/X16/9_X6/X14/X16/M8_s N_VDD_X6/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX6/X14/X16/M9 N_VDD_X6/X14/X16/M9_d N_X6/X14/19_X6/X14/X16/M9_g
+ N_X6/35_X6/X14/X16/M9_s N_VDD_X6/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/M0 N_GND_X7/M0_d N_X7/39_X7/M0_g N_X7/40_X7/M0_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/M1 N_X7/41_X7/M1_d N_X7/32_X7/M1_g N_GND_X7/M1_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12
mX7/M2 N_X7/42_X7/M2_d N_X7/31_X7/M2_g N_X7/41_X7/M2_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX7/M3 N_X7/43_X7/M3_d N_X7/30_X7/M3_g N_X7/42_X7/M3_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12
mX7/M4 N_X7/39_X7/M4_d N_X7/35_X7/M4_g N_X7/43_X7/M4_s N_GND_X0/X10/M0_b n
+ L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12
mX7/M5 N_VDD_X7/M5_d N_X7/39_X7/M5_g N_X7/40_X7/M5_s N_VDD_X7/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/M6 N_X7/39_X7/M6_d N_X7/32_X7/M6_g N_VDD_X7/M6_s N_VDD_X7/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX7/M7 N_VDD_X7/M7_d N_X7/31_X7/M7_g N_X7/39_X7/M7_s N_VDD_X7/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX7/M8 N_X7/39_X7/M8_d N_X7/30_X7/M8_g N_VDD_X7/M8_s N_VDD_X7/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12
mX7/M9 N_VDD_X7/M9_d N_X7/35_X7/M9_g N_X7/39_X7/M9_s N_VDD_X7/M5_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12
mX7/X10/M0 N_GND_X7/X10/M0_d N_9_X7/X10/M0_g N_51_X7/X10/M0_s N_GND_X0/X10/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X10/M1 N_X7/X10/10_X7/X10/M1_d N_C0_X7/X10/M1_g N_9_X7/X10/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X10/M2 N_GND_X7/X10/M2_d N_X7/40_X7/X10/M2_g N_X7/X10/10_X7/X10/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X10/M3 N_X7/X10/11_X7/X10/M3_d N_X7/39_X7/X10/M3_g N_GND_X7/X10/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X10/M4 N_9_X7/X10/M4_d N_X7/34_X7/X10/M4_g N_X7/X10/11_X7/X10/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X10/M5 N_X7/X10/9_X7/X10/M5_d N_X7/39_X7/X10/M5_g N_VDD_X7/X10/M5_s
+ N_VDD_X7/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX7/X10/M6 N_9_X7/X10/M6_d N_C0_X7/X10/M6_g N_X7/X10/9_X7/X10/M6_s
+ N_VDD_X7/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X10/M7 N_X7/X10/9_X7/X10/M7_d N_X7/40_X7/X10/M7_g N_9_X7/X10/M7_s
+ N_VDD_X7/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X10/M8 N_VDD_X7/X10/M8_d N_X7/34_X7/X10/M8_g N_X7/X10/9_X7/X10/M8_s
+ N_VDD_X7/X10/M5_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X10/M9 N_VDD_X7/X10/M9_d N_9_X7/X10/M9_g N_51_X7/X10/M9_s N_VDD_X7/X10/M5_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X11/M0 N_GND_X7/X11/M0_d N_X7/X11/14_X7/X11/M0_g N_X7/X11/16_X7/X11/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X11/M1 N_GND_X7/X11/M1_d N_X7/X11/13_X7/X11/M1_g N_X7/X11/14_X7/X11/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X11/M2 N_X7/X11/20_X7/X11/M2_d N_B2_X7/X11/M2_g N_GND_X7/X11/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X11/M3 N_X7/X11/14_X7/X11/M3_d N_A2_X7/X11/M3_g N_X7/X11/20_X7/X11/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X11/M4 N_GND_X7/X11/M4_d N_X7/X11/13_X7/X11/M4_g N_X7/X11/17_X7/X11/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X11/M5 N_X7/X11/13_X7/X11/M5_d N_B2_X7/X11/M5_g N_GND_X7/X11/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X11/M6 N_GND_X7/X11/M6_d N_A2_X7/X11/M6_g N_X7/X11/13_X7/X11/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X11/M7 N_X7/X11/15_X7/X11/M7_d N_X7/X11/13_X7/X11/M7_g
+ N_X7/X11/14_X7/X11/M7_s N_VDD_X7/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX7/X11/M8 N_VDD_X7/X11/M8_d N_B2_X7/X11/M8_g N_X7/X11/15_X7/X11/M8_s
+ N_VDD_X7/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X11/M9 N_X7/X11/15_X7/X11/M9_d N_A2_X7/X11/M9_g N_VDD_X7/X11/M9_s
+ N_VDD_X7/X11/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X11/M10 N_VDD_X7/X11/M10_d N_X7/X11/14_X7/X11/M10_g N_X7/X11/16_X7/X11/M10_s
+ N_VDD_X7/X11/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X11/M11 N_X7/X11/21_X7/X11/M11_d N_B2_X7/X11/M11_g N_VDD_X7/X11/M11_s
+ N_VDD_X7/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX7/X11/M12 N_X7/X11/13_X7/X11/M12_d N_A2_X7/X11/M12_g N_X7/X11/21_X7/X11/M12_s
+ N_VDD_X7/X11/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X11/M13 N_VDD_X7/X11/M13_d N_X7/X11/13_X7/X11/M13_g N_X7/X11/17_X7/X11/M13_s
+ N_VDD_X7/X11/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X11/X14/M0 N_GND_X7/X11/X14/M0_d N_X7/X11/18_X7/X11/X14/M0_g
+ N_SUM2_X7/X11/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X11/X14/M1 N_X7/X11/X14/10_X7/X11/X14/M1_d N_X7/30_X7/X11/X14/M1_g
+ N_X7/X11/18_X7/X11/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X11/X14/M2 N_GND_X7/X11/X14/M2_d N_X7/27_X7/X11/X14/M2_g
+ N_X7/X11/X14/10_X7/X11/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X11/X14/M3 N_X7/X11/X14/11_X7/X11/X14/M3_d N_X7/X11/16_X7/X11/X14/M3_g
+ N_GND_X7/X11/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X11/X14/M4 N_X7/X11/18_X7/X11/X14/M4_d N_X7/36_X7/X11/X14/M4_g
+ N_X7/X11/X14/11_X7/X11/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X11/X14/M5 N_X7/X11/X14/9_X7/X11/X14/M5_d N_X7/X11/16_X7/X11/X14/M5_g
+ N_VDD_X7/X11/X14/M5_s N_VDD_X7/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X11/X14/M6 N_X7/X11/18_X7/X11/X14/M6_d N_X7/30_X7/X11/X14/M6_g
+ N_X7/X11/X14/9_X7/X11/X14/M6_s N_VDD_X7/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X14/M7 N_X7/X11/X14/9_X7/X11/X14/M7_d N_X7/27_X7/X11/X14/M7_g
+ N_X7/X11/18_X7/X11/X14/M7_s N_VDD_X7/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X14/M8 N_VDD_X7/X11/X14/M8_d N_X7/36_X7/X11/X14/M8_g
+ N_X7/X11/X14/9_X7/X11/X14/M8_s N_VDD_X7/X11/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X11/X14/M9 N_VDD_X7/X11/X14/M9_d N_X7/X11/18_X7/X11/X14/M9_g
+ N_SUM2_X7/X11/X14/M9_s N_VDD_X7/X11/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X11/X15/M0 N_GND_X7/X11/X15/M0_d N_X7/29_X7/X11/X15/M0_g
+ N_X7/38_X7/X11/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X11/X15/M1 N_X7/X11/X15/10_X7/X11/X15/M1_d N_X7/X11/17_X7/X11/X15/M1_g
+ N_X7/29_X7/X11/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX7/X11/X15/M2 N_GND_X7/X11/X15/M2_d N_X7/36_X7/X11/X15/M2_g
+ N_X7/X11/X15/10_X7/X11/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X11/X15/M3 N_X7/X11/X15/11_X7/X11/X15/M3_d N_B2_X7/X11/X15/M3_g
+ N_GND_X7/X11/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X11/X15/M4 N_X7/29_X7/X11/X15/M4_d N_A2_X7/X11/X15/M4_g
+ N_X7/X11/X15/11_X7/X11/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X11/X15/M5 N_X7/X11/X15/9_X7/X11/X15/M5_d N_B2_X7/X11/X15/M5_g
+ N_VDD_X7/X11/X15/M5_s N_VDD_X7/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X11/X15/M6 N_X7/29_X7/X11/X15/M6_d N_X7/X11/17_X7/X11/X15/M6_g
+ N_X7/X11/X15/9_X7/X11/X15/M6_s N_VDD_X7/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X15/M7 N_X7/X11/X15/9_X7/X11/X15/M7_d N_X7/36_X7/X11/X15/M7_g
+ N_X7/29_X7/X11/X15/M7_s N_VDD_X7/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X15/M8 N_VDD_X7/X11/X15/M8_d N_A2_X7/X11/X15/M8_g
+ N_X7/X11/X15/9_X7/X11/X15/M8_s N_VDD_X7/X11/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X11/X15/M9 N_VDD_X7/X11/X15/M9_d N_X7/29_X7/X11/X15/M9_g
+ N_X7/38_X7/X11/X15/M9_s N_VDD_X7/X11/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X11/X16/M0 N_GND_X7/X11/X16/M0_d N_X7/X11/19_X7/X11/X16/M0_g
+ N_X7/30_X7/X11/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X11/X16/M1 N_X7/X11/X16/10_X7/X11/X16/M1_d N_A2N_X7/X11/X16/M1_g
+ N_X7/X11/19_X7/X11/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X11/X16/M2 N_GND_X7/X11/X16/M2_d N_B2_X7/X11/X16/M2_g
+ N_X7/X11/X16/10_X7/X11/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X11/X16/M3 N_X7/X11/X16/11_X7/X11/X16/M3_d N_B2N_X7/X11/X16/M3_g
+ N_GND_X7/X11/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X11/X16/M4 N_X7/X11/19_X7/X11/X16/M4_d N_A2_X7/X11/X16/M4_g
+ N_X7/X11/X16/11_X7/X11/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X11/X16/M5 N_X7/X11/X16/9_X7/X11/X16/M5_d N_B2N_X7/X11/X16/M5_g
+ N_VDD_X7/X11/X16/M5_s N_VDD_X7/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X11/X16/M6 N_X7/X11/19_X7/X11/X16/M6_d N_A2N_X7/X11/X16/M6_g
+ N_X7/X11/X16/9_X7/X11/X16/M6_s N_VDD_X7/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X16/M7 N_X7/X11/X16/9_X7/X11/X16/M7_d N_B2_X7/X11/X16/M7_g
+ N_X7/X11/19_X7/X11/X16/M7_s N_VDD_X7/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X11/X16/M8 N_VDD_X7/X11/X16/M8_d N_A2_X7/X11/X16/M8_g
+ N_X7/X11/X16/9_X7/X11/X16/M8_s N_VDD_X7/X11/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X11/X16/M9 N_VDD_X7/X11/X16/M9_d N_X7/X11/19_X7/X11/X16/M9_g
+ N_X7/30_X7/X11/X16/M9_s N_VDD_X7/X11/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X12/M0 N_GND_X7/X12/M0_d N_X7/X12/14_X7/X12/M0_g N_X7/X12/16_X7/X12/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X12/M1 N_GND_X7/X12/M1_d N_X7/X12/13_X7/X12/M1_g N_X7/X12/14_X7/X12/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X12/M2 N_X7/X12/20_X7/X12/M2_d N_B1_X7/X12/M2_g N_GND_X7/X12/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X12/M3 N_X7/X12/14_X7/X12/M3_d N_A1_X7/X12/M3_g N_X7/X12/20_X7/X12/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X12/M4 N_GND_X7/X12/M4_d N_X7/X12/13_X7/X12/M4_g N_X7/X12/17_X7/X12/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X12/M5 N_X7/X12/13_X7/X12/M5_d N_B1_X7/X12/M5_g N_GND_X7/X12/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X12/M6 N_GND_X7/X12/M6_d N_A1_X7/X12/M6_g N_X7/X12/13_X7/X12/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X12/M7 N_X7/X12/15_X7/X12/M7_d N_X7/X12/13_X7/X12/M7_g
+ N_X7/X12/14_X7/X12/M7_s N_VDD_X7/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX7/X12/M8 N_VDD_X7/X12/M8_d N_B1_X7/X12/M8_g N_X7/X12/15_X7/X12/M8_s
+ N_VDD_X7/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X12/M9 N_X7/X12/15_X7/X12/M9_d N_A1_X7/X12/M9_g N_VDD_X7/X12/M9_s
+ N_VDD_X7/X12/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X12/M10 N_VDD_X7/X12/M10_d N_X7/X12/14_X7/X12/M10_g N_X7/X12/16_X7/X12/M10_s
+ N_VDD_X7/X12/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X12/M11 N_X7/X12/21_X7/X12/M11_d N_B1_X7/X12/M11_g N_VDD_X7/X12/M11_s
+ N_VDD_X7/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX7/X12/M12 N_X7/X12/13_X7/X12/M12_d N_A1_X7/X12/M12_g N_X7/X12/21_X7/X12/M12_s
+ N_VDD_X7/X12/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X12/M13 N_VDD_X7/X12/M13_d N_X7/X12/13_X7/X12/M13_g N_X7/X12/17_X7/X12/M13_s
+ N_VDD_X7/X12/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X12/X14/M0 N_GND_X7/X12/X14/M0_d N_X7/X12/18_X7/X12/X14/M0_g
+ N_SUM1_X7/X12/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X12/X14/M1 N_X7/X12/X14/10_X7/X12/X14/M1_d N_X7/31_X7/X12/X14/M1_g
+ N_X7/X12/18_X7/X12/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X12/X14/M2 N_GND_X7/X12/X14/M2_d N_X7/28_X7/X12/X14/M2_g
+ N_X7/X12/X14/10_X7/X12/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X12/X14/M3 N_X7/X12/X14/11_X7/X12/X14/M3_d N_X7/X12/16_X7/X12/X14/M3_g
+ N_GND_X7/X12/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X12/X14/M4 N_X7/X12/18_X7/X12/X14/M4_d N_X7/37_X7/X12/X14/M4_g
+ N_X7/X12/X14/11_X7/X12/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X12/X14/M5 N_X7/X12/X14/9_X7/X12/X14/M5_d N_X7/X12/16_X7/X12/X14/M5_g
+ N_VDD_X7/X12/X14/M5_s N_VDD_X7/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X12/X14/M6 N_X7/X12/18_X7/X12/X14/M6_d N_X7/31_X7/X12/X14/M6_g
+ N_X7/X12/X14/9_X7/X12/X14/M6_s N_VDD_X7/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X14/M7 N_X7/X12/X14/9_X7/X12/X14/M7_d N_X7/28_X7/X12/X14/M7_g
+ N_X7/X12/18_X7/X12/X14/M7_s N_VDD_X7/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X14/M8 N_VDD_X7/X12/X14/M8_d N_X7/37_X7/X12/X14/M8_g
+ N_X7/X12/X14/9_X7/X12/X14/M8_s N_VDD_X7/X12/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X12/X14/M9 N_VDD_X7/X12/X14/M9_d N_X7/X12/18_X7/X12/X14/M9_g
+ N_SUM1_X7/X12/X14/M9_s N_VDD_X7/X12/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X12/X15/M0 N_GND_X7/X12/X15/M0_d N_X7/27_X7/X12/X15/M0_g
+ N_X7/36_X7/X12/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X12/X15/M1 N_X7/X12/X15/10_X7/X12/X15/M1_d N_X7/X12/17_X7/X12/X15/M1_g
+ N_X7/27_X7/X12/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX7/X12/X15/M2 N_GND_X7/X12/X15/M2_d N_X7/37_X7/X12/X15/M2_g
+ N_X7/X12/X15/10_X7/X12/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X12/X15/M3 N_X7/X12/X15/11_X7/X12/X15/M3_d N_B1_X7/X12/X15/M3_g
+ N_GND_X7/X12/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X12/X15/M4 N_X7/27_X7/X12/X15/M4_d N_A1_X7/X12/X15/M4_g
+ N_X7/X12/X15/11_X7/X12/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X12/X15/M5 N_X7/X12/X15/9_X7/X12/X15/M5_d N_B1_X7/X12/X15/M5_g
+ N_VDD_X7/X12/X15/M5_s N_VDD_X7/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X12/X15/M6 N_X7/27_X7/X12/X15/M6_d N_X7/X12/17_X7/X12/X15/M6_g
+ N_X7/X12/X15/9_X7/X12/X15/M6_s N_VDD_X7/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X15/M7 N_X7/X12/X15/9_X7/X12/X15/M7_d N_X7/37_X7/X12/X15/M7_g
+ N_X7/27_X7/X12/X15/M7_s N_VDD_X7/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X15/M8 N_VDD_X7/X12/X15/M8_d N_A1_X7/X12/X15/M8_g
+ N_X7/X12/X15/9_X7/X12/X15/M8_s N_VDD_X7/X12/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X12/X15/M9 N_VDD_X7/X12/X15/M9_d N_X7/27_X7/X12/X15/M9_g
+ N_X7/36_X7/X12/X15/M9_s N_VDD_X7/X12/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X12/X16/M0 N_GND_X7/X12/X16/M0_d N_X7/X12/19_X7/X12/X16/M0_g
+ N_X7/31_X7/X12/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X12/X16/M1 N_X7/X12/X16/10_X7/X12/X16/M1_d N_A1N_X7/X12/X16/M1_g
+ N_X7/X12/19_X7/X12/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X12/X16/M2 N_GND_X7/X12/X16/M2_d N_B1_X7/X12/X16/M2_g
+ N_X7/X12/X16/10_X7/X12/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X12/X16/M3 N_X7/X12/X16/11_X7/X12/X16/M3_d N_B1N_X7/X12/X16/M3_g
+ N_GND_X7/X12/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X12/X16/M4 N_X7/X12/19_X7/X12/X16/M4_d N_A1_X7/X12/X16/M4_g
+ N_X7/X12/X16/11_X7/X12/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X12/X16/M5 N_X7/X12/X16/9_X7/X12/X16/M5_d N_B1N_X7/X12/X16/M5_g
+ N_VDD_X7/X12/X16/M5_s N_VDD_X7/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X12/X16/M6 N_X7/X12/19_X7/X12/X16/M6_d N_A1N_X7/X12/X16/M6_g
+ N_X7/X12/X16/9_X7/X12/X16/M6_s N_VDD_X7/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X16/M7 N_X7/X12/X16/9_X7/X12/X16/M7_d N_B1_X7/X12/X16/M7_g
+ N_X7/X12/19_X7/X12/X16/M7_s N_VDD_X7/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X12/X16/M8 N_VDD_X7/X12/X16/M8_d N_A1_X7/X12/X16/M8_g
+ N_X7/X12/X16/9_X7/X12/X16/M8_s N_VDD_X7/X12/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X12/X16/M9 N_VDD_X7/X12/X16/M9_d N_X7/X12/19_X7/X12/X16/M9_g
+ N_X7/31_X7/X12/X16/M9_s N_VDD_X7/X12/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X13/M0 N_GND_X7/X13/M0_d N_X7/X13/14_X7/X13/M0_g N_X7/X13/16_X7/X13/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X13/M1 N_GND_X7/X13/M1_d N_X7/X13/13_X7/X13/M1_g N_X7/X13/14_X7/X13/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X13/M2 N_X7/X13/20_X7/X13/M2_d N_B0_X7/X13/M2_g N_GND_X7/X13/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X13/M3 N_X7/X13/14_X7/X13/M3_d N_A0_X7/X13/M3_g N_X7/X13/20_X7/X13/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X13/M4 N_GND_X7/X13/M4_d N_X7/X13/13_X7/X13/M4_g N_X7/X13/17_X7/X13/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X13/M5 N_X7/X13/13_X7/X13/M5_d N_B0_X7/X13/M5_g N_GND_X7/X13/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X13/M6 N_GND_X7/X13/M6_d N_A0_X7/X13/M6_g N_X7/X13/13_X7/X13/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X13/M7 N_X7/X13/15_X7/X13/M7_d N_X7/X13/13_X7/X13/M7_g
+ N_X7/X13/14_X7/X13/M7_s N_VDD_X7/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX7/X13/M8 N_VDD_X7/X13/M8_d N_B0_X7/X13/M8_g N_X7/X13/15_X7/X13/M8_s
+ N_VDD_X7/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X13/M9 N_X7/X13/15_X7/X13/M9_d N_A0_X7/X13/M9_g N_VDD_X7/X13/M9_s
+ N_VDD_X7/X13/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X13/M10 N_VDD_X7/X13/M10_d N_X7/X13/14_X7/X13/M10_g N_X7/X13/16_X7/X13/M10_s
+ N_VDD_X7/X13/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X13/M11 N_X7/X13/21_X7/X13/M11_d N_B0_X7/X13/M11_g N_VDD_X7/X13/M11_s
+ N_VDD_X7/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX7/X13/M12 N_X7/X13/13_X7/X13/M12_d N_A0_X7/X13/M12_g N_X7/X13/21_X7/X13/M12_s
+ N_VDD_X7/X13/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X13/M13 N_VDD_X7/X13/M13_d N_X7/X13/13_X7/X13/M13_g N_X7/X13/17_X7/X13/M13_s
+ N_VDD_X7/X13/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X13/X14/M0 N_GND_X7/X13/X14/M0_d N_X7/X13/18_X7/X13/X14/M0_g
+ N_SUM0_X7/X13/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X13/X14/M1 N_X7/X13/X14/10_X7/X13/X14/M1_d N_X7/32_X7/X13/X14/M1_g
+ N_X7/X13/18_X7/X13/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X13/X14/M2 N_GND_X7/X13/X14/M2_d N_C0N_X7/X13/X14/M2_g
+ N_X7/X13/X14/10_X7/X13/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X13/X14/M3 N_X7/X13/X14/11_X7/X13/X14/M3_d N_X7/X13/16_X7/X13/X14/M3_g
+ N_GND_X7/X13/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X13/X14/M4 N_X7/X13/18_X7/X13/X14/M4_d N_C0_X7/X13/X14/M4_g
+ N_X7/X13/X14/11_X7/X13/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X13/X14/M5 N_X7/X13/X14/9_X7/X13/X14/M5_d N_X7/X13/16_X7/X13/X14/M5_g
+ N_VDD_X7/X13/X14/M5_s N_VDD_X7/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X13/X14/M6 N_X7/X13/18_X7/X13/X14/M6_d N_X7/32_X7/X13/X14/M6_g
+ N_X7/X13/X14/9_X7/X13/X14/M6_s N_VDD_X7/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X14/M7 N_X7/X13/X14/9_X7/X13/X14/M7_d N_C0N_X7/X13/X14/M7_g
+ N_X7/X13/18_X7/X13/X14/M7_s N_VDD_X7/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X14/M8 N_VDD_X7/X13/X14/M8_d N_C0_X7/X13/X14/M8_g
+ N_X7/X13/X14/9_X7/X13/X14/M8_s N_VDD_X7/X13/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X13/X14/M9 N_VDD_X7/X13/X14/M9_d N_X7/X13/18_X7/X13/X14/M9_g
+ N_SUM0_X7/X13/X14/M9_s N_VDD_X7/X13/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X13/X15/M0 N_GND_X7/X13/X15/M0_d N_X7/28_X7/X13/X15/M0_g
+ N_X7/37_X7/X13/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X13/X15/M1 N_X7/X13/X15/10_X7/X13/X15/M1_d N_X7/X13/17_X7/X13/X15/M1_g
+ N_X7/28_X7/X13/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX7/X13/X15/M2 N_GND_X7/X13/X15/M2_d N_C0_X7/X13/X15/M2_g
+ N_X7/X13/X15/10_X7/X13/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X13/X15/M3 N_X7/X13/X15/11_X7/X13/X15/M3_d N_B0_X7/X13/X15/M3_g
+ N_GND_X7/X13/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X13/X15/M4 N_X7/28_X7/X13/X15/M4_d N_A0_X7/X13/X15/M4_g
+ N_X7/X13/X15/11_X7/X13/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X13/X15/M5 N_X7/X13/X15/9_X7/X13/X15/M5_d N_B0_X7/X13/X15/M5_g
+ N_VDD_X7/X13/X15/M5_s N_VDD_X7/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X13/X15/M6 N_X7/28_X7/X13/X15/M6_d N_X7/X13/17_X7/X13/X15/M6_g
+ N_X7/X13/X15/9_X7/X13/X15/M6_s N_VDD_X7/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X15/M7 N_X7/X13/X15/9_X7/X13/X15/M7_d N_C0_X7/X13/X15/M7_g
+ N_X7/28_X7/X13/X15/M7_s N_VDD_X7/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X15/M8 N_VDD_X7/X13/X15/M8_d N_A0_X7/X13/X15/M8_g
+ N_X7/X13/X15/9_X7/X13/X15/M8_s N_VDD_X7/X13/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X13/X15/M9 N_VDD_X7/X13/X15/M9_d N_X7/28_X7/X13/X15/M9_g
+ N_X7/37_X7/X13/X15/M9_s N_VDD_X7/X13/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X13/X16/M0 N_GND_X7/X13/X16/M0_d N_X7/X13/19_X7/X13/X16/M0_g
+ N_X7/32_X7/X13/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X13/X16/M1 N_X7/X13/X16/10_X7/X13/X16/M1_d N_A0N_X7/X13/X16/M1_g
+ N_X7/X13/19_X7/X13/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X13/X16/M2 N_GND_X7/X13/X16/M2_d N_B0_X7/X13/X16/M2_g
+ N_X7/X13/X16/10_X7/X13/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X13/X16/M3 N_X7/X13/X16/11_X7/X13/X16/M3_d N_B0N_X7/X13/X16/M3_g
+ N_GND_X7/X13/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X13/X16/M4 N_X7/X13/19_X7/X13/X16/M4_d N_A0_X7/X13/X16/M4_g
+ N_X7/X13/X16/11_X7/X13/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X13/X16/M5 N_X7/X13/X16/9_X7/X13/X16/M5_d N_B0N_X7/X13/X16/M5_g
+ N_VDD_X7/X13/X16/M5_s N_VDD_X7/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X13/X16/M6 N_X7/X13/19_X7/X13/X16/M6_d N_A0N_X7/X13/X16/M6_g
+ N_X7/X13/X16/9_X7/X13/X16/M6_s N_VDD_X7/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X16/M7 N_X7/X13/X16/9_X7/X13/X16/M7_d N_B0_X7/X13/X16/M7_g
+ N_X7/X13/19_X7/X13/X16/M7_s N_VDD_X7/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X13/X16/M8 N_VDD_X7/X13/X16/M8_d N_A0_X7/X13/X16/M8_g
+ N_X7/X13/X16/9_X7/X13/X16/M8_s N_VDD_X7/X13/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X13/X16/M9 N_VDD_X7/X13/X16/M9_d N_X7/X13/19_X7/X13/X16/M9_g
+ N_X7/32_X7/X13/X16/M9_s N_VDD_X7/X13/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X14/M0 N_GND_X7/X14/M0_d N_X7/X14/14_X7/X14/M0_g N_X7/X14/16_X7/X14/M0_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X14/M1 N_GND_X7/X14/M1_d N_X7/X14/13_X7/X14/M1_g N_X7/X14/14_X7/X14/M1_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X14/M2 N_X7/X14/20_X7/X14/M2_d N_B3_X7/X14/M2_g N_GND_X7/X14/M2_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13
mX7/X14/M3 N_X7/X14/14_X7/X14/M3_d N_A3_X7/X14/M3_g N_X7/X14/20_X7/X14/M3_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X14/M4 N_GND_X7/X14/M4_d N_X7/X14/13_X7/X14/M4_g N_X7/X14/17_X7/X14/M4_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X14/M5 N_X7/X14/13_X7/X14/M5_d N_B3_X7/X14/M5_g N_GND_X7/X14/M5_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13
mX7/X14/M6 N_GND_X7/X14/M6_d N_A3_X7/X14/M6_g N_X7/X14/13_X7/X14/M6_s
+ N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13
mX7/X14/M7 N_X7/X14/15_X7/X14/M7_d N_X7/X14/13_X7/X14/M7_g
+ N_X7/X14/14_X7/X14/M7_s N_VDD_X7/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12
+ AS=2.3328e-12
mX7/X14/M8 N_VDD_X7/X14/M8_d N_B3_X7/X14/M8_g N_X7/X14/15_X7/X14/M8_s
+ N_VDD_X7/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12
mX7/X14/M9 N_X7/X14/15_X7/X14/M9_d N_A3_X7/X14/M9_g N_VDD_X7/X14/M9_s
+ N_VDD_X7/X14/M7_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X14/M10 N_VDD_X7/X14/M10_d N_X7/X14/14_X7/X14/M10_g N_X7/X14/16_X7/X14/M10_s
+ N_VDD_X7/X14/M7_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X14/M11 N_X7/X14/21_X7/X14/M11_d N_B3_X7/X14/M11_g N_VDD_X7/X14/M11_s
+ N_VDD_X7/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12
mX7/X14/M12 N_X7/X14/13_X7/X14/M12_d N_A3_X7/X14/M12_g N_X7/X14/21_X7/X14/M12_s
+ N_VDD_X7/X14/M11_b p L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12
mX7/X14/M13 N_VDD_X7/X14/M13_d N_X7/X14/13_X7/X14/M13_g N_X7/X14/17_X7/X14/M13_s
+ N_VDD_X7/X14/M11_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X14/X14/M0 N_GND_X7/X14/X14/M0_d N_X7/X14/18_X7/X14/X14/M0_g
+ N_SUM3_X7/X14/X14/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X14/X14/M1 N_X7/X14/X14/10_X7/X14/X14/M1_d N_X7/35_X7/X14/X14/M1_g
+ N_X7/X14/18_X7/X14/X14/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X14/X14/M2 N_GND_X7/X14/X14/M2_d N_X7/29_X7/X14/X14/M2_g
+ N_X7/X14/X14/10_X7/X14/X14/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X14/X14/M3 N_X7/X14/X14/11_X7/X14/X14/M3_d N_X7/X14/16_X7/X14/X14/M3_g
+ N_GND_X7/X14/X14/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X14/X14/M4 N_X7/X14/18_X7/X14/X14/M4_d N_X7/38_X7/X14/X14/M4_g
+ N_X7/X14/X14/11_X7/X14/X14/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X14/X14/M5 N_X7/X14/X14/9_X7/X14/X14/M5_d N_X7/X14/16_X7/X14/X14/M5_g
+ N_VDD_X7/X14/X14/M5_s N_VDD_X7/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X14/X14/M6 N_X7/X14/18_X7/X14/X14/M6_d N_X7/35_X7/X14/X14/M6_g
+ N_X7/X14/X14/9_X7/X14/X14/M6_s N_VDD_X7/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X14/M7 N_X7/X14/X14/9_X7/X14/X14/M7_d N_X7/29_X7/X14/X14/M7_g
+ N_X7/X14/18_X7/X14/X14/M7_s N_VDD_X7/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X14/M8 N_VDD_X7/X14/X14/M8_d N_X7/38_X7/X14/X14/M8_g
+ N_X7/X14/X14/9_X7/X14/X14/M8_s N_VDD_X7/X14/X14/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X14/X14/M9 N_VDD_X7/X14/X14/M9_d N_X7/X14/18_X7/X14/X14/M9_g
+ N_SUM3_X7/X14/X14/M9_s N_VDD_X7/X14/X14/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X14/X15/M0 N_GND_X7/X14/X15/M0_d N_X7/33_X7/X14/X15/M0_g
+ N_X7/34_X7/X14/X15/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X14/X15/M1 N_X7/X14/X15/10_X7/X14/X15/M1_d N_X7/X14/17_X7/X14/X15/M1_g
+ N_X7/33_X7/X14/X15/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
mX7/X14/X15/M2 N_GND_X7/X14/X15/M2_d N_X7/38_X7/X14/X15/M2_g
+ N_X7/X14/X15/10_X7/X14/X15/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X14/X15/M3 N_X7/X14/X15/11_X7/X14/X15/M3_d N_B3_X7/X14/X15/M3_g
+ N_GND_X7/X14/X15/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X14/X15/M4 N_X7/33_X7/X14/X15/M4_d N_A3_X7/X14/X15/M4_g
+ N_X7/X14/X15/11_X7/X14/X15/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X14/X15/M5 N_X7/X14/X15/9_X7/X14/X15/M5_d N_B3_X7/X14/X15/M5_g
+ N_VDD_X7/X14/X15/M5_s N_VDD_X7/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X14/X15/M6 N_X7/33_X7/X14/X15/M6_d N_X7/X14/17_X7/X14/X15/M6_g
+ N_X7/X14/X15/9_X7/X14/X15/M6_s N_VDD_X7/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X15/M7 N_X7/X14/X15/9_X7/X14/X15/M7_d N_X7/38_X7/X14/X15/M7_g
+ N_X7/33_X7/X14/X15/M7_s N_VDD_X7/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X15/M8 N_VDD_X7/X14/X15/M8_d N_A3_X7/X14/X15/M8_g
+ N_X7/X14/X15/9_X7/X14/X15/M8_s N_VDD_X7/X14/X15/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X14/X15/M9 N_VDD_X7/X14/X15/M9_d N_X7/33_X7/X14/X15/M9_g
+ N_X7/34_X7/X14/X15/M9_s N_VDD_X7/X14/X15/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
mX7/X14/X16/M0 N_GND_X7/X14/X16/M0_d N_X7/X14/19_X7/X14/X16/M0_g
+ N_X7/35_X7/X14/X16/M0_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=4.374e-13
mX7/X14/X16/M1 N_X7/X14/X16/10_X7/X14/X16/M1_d N_A3N_X7/X14/X16/M1_g
+ N_X7/X14/19_X7/X14/X16/M1_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
mX7/X14/X16/M2 N_GND_X7/X14/X16/M2_d N_B3_X7/X14/X16/M2_g
+ N_X7/X14/X16/10_X7/X14/X16/M2_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
mX7/X14/X16/M3 N_X7/X14/X16/11_X7/X14/X16/M3_d N_B3N_X7/X14/X16/M3_g
+ N_GND_X7/X14/X16/M3_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
mX7/X14/X16/M4 N_X7/X14/19_X7/X14/X16/M4_d N_A3_X7/X14/X16/M4_g
+ N_X7/X14/X16/11_X7/X14/X16/M4_s N_GND_X0/X10/M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
mX7/X14/X16/M5 N_X7/X14/X16/9_X7/X14/X16/M5_d N_B3N_X7/X14/X16/M5_g
+ N_VDD_X7/X14/X16/M5_s N_VDD_X7/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
mX7/X14/X16/M6 N_X7/X14/19_X7/X14/X16/M6_d N_A3N_X7/X14/X16/M6_g
+ N_X7/X14/X16/9_X7/X14/X16/M6_s N_VDD_X7/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X16/M7 N_X7/X14/X16/9_X7/X14/X16/M7_d N_B3_X7/X14/X16/M7_g
+ N_X7/X14/19_X7/X14/X16/M7_s N_VDD_X7/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
mX7/X14/X16/M8 N_VDD_X7/X14/X16/M8_d N_A3_X7/X14/X16/M8_g
+ N_X7/X14/X16/9_X7/X14/X16/M8_s N_VDD_X7/X14/X16/M5_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
mX7/X14/X16/M9 N_VDD_X7/X14/X16/M9_d N_X7/X14/19_X7/X14/X16/M9_g
+ N_X7/35_X7/X14/X16/M9_s N_VDD_X7/X14/X16/M5_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
*
.include "thirty_two_bit_adder.pex.netlist.THIRTY_TWO_BIT_ADDER.pxi"
*
.ends
*
*
