* SPICE NETLIST
***************************************

.SUBCKT i VDD IN2 IN4 IN3 IN1 OUTN OUT GND
** N=11 EP=8 IP=0 FDC=10
* PORT VDD VDD -23500 1500 METAL2
* PORT IN2 IN2 -21000 30000 METAL1
* PORT IN2 IN2 151000 58000 METAL1
* PORT IN4 IN4 -21000 44000 METAL1
* PORT IN4 IN4 151000 30000 METAL1
* PORT IN3 IN3 -21000 58000 METAL1
* PORT IN3 IN3 151000 44000 METAL1
* PORT IN1 IN1 -21000 72000 METAL1
* PORT IN1 IN1 151000 72000 METAL1
* PORT OUTN OUTN 37000 -33000 METAL1
* PORT OUT OUT 79000 -33000 METAL1
* PORT GND GND 151000 10000 METAL1
M0 GND OUTN OUT GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=90000 $Y=-12000 $D=1
M1 10 IN4 OUTN GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=113000 $Y=29000 $D=1
M2 GND IN3 10 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=43000 $D=1
M3 11 IN2 GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=57000 $D=1
M4 OUTN IN1 11 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=113000 $Y=71000 $D=1
M5 9 IN2 VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=33000 $Y=29000 $D=0
M6 OUTN IN4 9 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=43000 $D=0
M7 9 IN3 OUTN VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=57000 $D=0
M8 VDD IN1 9 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=33000 $Y=71000 $D=0
M9 VDD OUTN OUT VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=49000 $Y=-12000 $D=0
.ENDS
***************************************
.SUBCKT full_adder COUTN CN COUT C VDD GND SUM B A P AN BN
** N=21 EP=12 IP=24 FDC=44
* PORT COUTN COUTN 269500 -18000 METAL2
* PORT CN CN 286500 207500 METAL2
* PORT COUT COUT 311500 -18000 METAL1
* PORT C C 403000 190000 METAL1
* PORT VDD VDD -493000 90500 METAL1
* PORT GND GND 648000 98500 METAL1
* PORT SUM SUM -493000 29500 METAL1
* PORT B B 648000 132500 METAL1
* PORT A A 648000 160500 METAL1
* PORT P P 560000 -18000 METAL1
* PORT AN AN 648000 118500 METAL1
* PORT BN BN 648000 146500 METAL1
M0 GND 14 16 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=-121000 $Y=75000 $D=1
M1 GND 13 14 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=-118000 $Y=119000 $D=1
M2 20 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=-118000 $Y=133000 $D=1
M3 14 A 20 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=-118000 $Y=147000 $D=1
M4 GND 13 17 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=81000 $Y=76500 $D=1
M5 13 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=92000 $Y=117500 $D=1
M6 GND A 13 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=92000 $Y=131500 $D=1
M7 15 13 14 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=-177000 $Y=119000 $D=0
M8 VDD B 15 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=-177000 $Y=133000 $D=0
M9 15 A VDD VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=-177000 $Y=147000 $D=0
M10 VDD 14 16 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-162000 $Y=75000 $D=0
M11 21 B VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=31000 $Y=117500 $D=0
M12 13 A 21 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=31000 $Y=131500 $D=0
M13 VDD 13 17 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=47000 $Y=76500 $D=0
X14 VDD 16 P CN C 18 SUM GND i $T=-438000 89000 0 0 $X=-464000 $Y=54000
X15 VDD B 17 C A COUTN COUT GND i $T=232500 85000 0 0 $X=206500 $Y=50000
X16 VDD BN AN B A 19 P GND i $T=481000 88500 0 0 $X=455000 $Y=53500
.ENDS
***************************************
.SUBCKT four_bit_adder VDD COUTN C0N C0 GND SUM2 SUM1 SUM0 SUM3 COUT A2N B2 B2N A2 A1N B1 B1N A1 A0N B0
+ B0N A0 A3N B3 B3N A3
** N=43 EP=26 IP=56 FDC=196
* PORT VDD VDD 282000 508000 METAL2
* PORT VDD VDD 302500 -792000 METAL2
* PORT COUTN COUTN 979000 -798000 METAL2
* PORT C0N C0N 1134000 527000 METAL2
* PORT C0 C0 1250500 527000 METAL1
* PORT GND GND 1811000 519500 METAL2
* PORT GND GND 1817000 -786000 METAL2
* PORT SUM2 SUM2 218500 -224000 METAL1
* PORT SUM1 SUM1 220000 61500 METAL1
* PORT SUM0 SUM0 222000 333500 METAL1
* PORT SUM3 SUM3 224000 -509000 METAL1
* PORT COUT COUT 1021000 -798000 METAL1
* PORT A2N A2N 1894500 -135000 METAL1
* PORT B2 B2 1894500 -121000 METAL1
* PORT B2N B2N 1894500 -107000 METAL1
* PORT A2 A2 1894500 -93000 METAL1
* PORT A1N A1N 1896000 150500 METAL1
* PORT B1 B1 1896000 164500 METAL1
* PORT B1N B1N 1896000 178500 METAL1
* PORT A1 A1 1896000 192500 METAL1
* PORT A0N A0N 1898000 422500 METAL1
* PORT B0 B0 1898000 436500 METAL1
* PORT B0N B0N 1898000 450500 METAL1
* PORT A0 A0 1898000 464500 METAL1
* PORT A3N A3N 1900000 -420000 METAL1
* PORT B3 B3 1900000 -406000 METAL1
* PORT B3N B3N 1900000 -392000 METAL1
* PORT A3 A3 1900000 -378000 METAL1
M0 GND 39 40 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=1307500 $Y=-714000 $D=1
M1 41 32 GND GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12 $X=1310500 $Y=-675000 $D=1
M2 42 31 41 GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12 $X=1310500 $Y=-661000 $D=1
M3 43 30 42 GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12 $X=1310500 $Y=-647000 $D=1
M4 39 35 43 GND N L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12 $X=1310500 $Y=-633000 $D=1
M5 VDD 39 40 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=1266500 $Y=-714000 $D=0
M6 39 32 VDD VDD P L=1.8e-07 W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12 $X=1268500 $Y=-675000 $D=0
M7 VDD 31 39 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12 $X=1268500 $Y=-661000 $D=0
M8 39 30 VDD VDD P L=1.8e-07 W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12 $X=1268500 $Y=-631000 $D=0
M9 VDD 35 39 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12 $X=1268500 $Y=-617000 $D=0
X10 VDD 39 C0 40 34 COUTN COUT GND i $T=942000 -686000 0 0 $X=916000 $Y=-721000
X11 29 27 38 36 VDD GND SUM2 B2 A2 30 A2N B2N full_adder $T=844000 -253500 0 0 $X=349000 $Y=-273500
X12 27 28 36 37 VDD GND SUM1 B1 A1 31 A1N B1N full_adder $T=845500 32000 0 0 $X=350500 $Y=12000
X13 28 C0N 37 C0 VDD GND SUM0 B0 A0 32 A0N B0N full_adder $T=847500 304000 0 0 $X=352500 $Y=284000
X14 33 29 34 38 VDD GND SUM3 B3 A3 35 A3N B3N full_adder $T=849500 -538500 0 0 $X=354500 $Y=-558500
.ENDS
***************************************
.SUBCKT thirty_two_bit_adder VDD COUT31N C0N GND SUM30 SUM26 SUM22 SUM29 SUM25 SUM21 SUM28 SUM24 SUM20 SUM31 SUM27 SUM23 SUM14 SUM10 SUM18 SUM6
+ SUM13 SUM9 SUM17 SUM5 SUM12 SUM8 SUM16 SUM4 SUM15 SUM11 SUM19 SUM7 SUM2 SUM1 SUM0 SUM3 COUT31 C0 A30N B30
+ B30N A30 A26N B26 B26N A26 A22N B22 B22N A22 A29N B29 B29N A29 A25N B25 B25N A25 A21N B21
+ B21N A21 A28N B28 B28N A28 A24N B24 B24N A24 A20N B20 B20N A20 A31N B31 B31N A31 A27N B27
+ B27N A27 A23N B23 B23N A23 A14N B14 B14N A14 A10N B10 B10N A10 A18N B18 B18N A18 A6N B6
+ B6N A6 A13N B13 B13N A13 A9N B9 B9N A9 A17N B17 B17N A17 A5N B5 B5N A5 A12N B12
+ B12N A12 A8N B8 B8N A8 A16N B16 B16N A16 A4N B4 B4N A4 A15N B15 B15N A15 A11N B11
+ B11N A11 A19N B19 B19N A19 A7N B7 B7N A7 A2N B2 B2N A2 A1N B1 B1N A1 A0N B0
+ B0N A0 A3N B3 B3N A3
** N=180 EP=166 IP=208 FDC=1568
* PORT VDD VDD 528000 1508000 METAL2
* PORT COUT31N COUT31N 1211500 -9878000 METAL2
* PORT C0N C0N 1380000 1513000 METAL2
* PORT GND GND 2057000 1513000 METAL2
* PORT SUM30 SUM30 425000 -9254500 METAL1
* PORT SUM26 SUM26 425000 -7839000 METAL1
* PORT SUM22 SUM22 425500 -6393500 METAL1
* PORT SUM29 SUM29 426500 -8969000 METAL1
* PORT SUM25 SUM25 426500 -7553500 METAL1
* PORT SUM21 SUM21 427000 -6108000 METAL1
* PORT SUM28 SUM28 428500 -8697000 METAL1
* PORT SUM24 SUM24 428500 -7281500 METAL1
* PORT SUM20 SUM20 429000 -5836000 METAL1
* PORT SUM31 SUM31 430500 -9539500 METAL1
* PORT SUM27 SUM27 430500 -8124000 METAL1
* PORT SUM23 SUM23 431000 -6678500 METAL1
* PORT SUM14 SUM14 431500 -3526500 METAL1
* PORT SUM10 SUM10 431500 -2111000 METAL1
* PORT SUM18 SUM18 432000 -4988500 METAL1
* PORT SUM6 SUM6 432000 -665500 METAL1
* PORT SUM13 SUM13 433000 -3241000 METAL1
* PORT SUM9 SUM9 433000 -1825500 METAL1
* PORT SUM17 SUM17 433500 -4703000 METAL1
* PORT SUM5 SUM5 433500 -380000 METAL1
* PORT SUM12 SUM12 435000 -2969000 METAL1
* PORT SUM8 SUM8 435000 -1553500 METAL1
* PORT SUM16 SUM16 435500 -4431000 METAL1
* PORT SUM4 SUM4 435500 -108000 METAL1
* PORT SUM15 SUM15 437000 -3811500 METAL1
* PORT SUM11 SUM11 437000 -2396000 METAL1
* PORT SUM19 SUM19 437500 -5273500 METAL1
* PORT SUM7 SUM7 437500 -950500 METAL1
* PORT SUM2 SUM2 438500 739500 METAL1
* PORT SUM1 SUM1 440000 1025000 METAL1
* PORT SUM0 SUM0 442000 1297000 METAL1
* PORT SUM3 SUM3 444000 454500 METAL1
* PORT COUT31 COUT31 1253500 -9878000 METAL1
* PORT C0 C0 1496500 1513000 METAL1
* PORT A30N A30N 2154500 -9165500 METAL1
* PORT B30 B30 2154500 -9151500 METAL1
* PORT B30N B30N 2154500 -9137500 METAL1
* PORT A30 A30 2154500 -9123500 METAL1
* PORT A26N A26N 2154500 -7750000 METAL1
* PORT B26 B26 2154500 -7736000 METAL1
* PORT B26N B26N 2154500 -7722000 METAL1
* PORT A26 A26 2154500 -7708000 METAL1
* PORT A22N A22N 2155000 -6304500 METAL1
* PORT B22 B22 2155000 -6290500 METAL1
* PORT B22N B22N 2155000 -6276500 METAL1
* PORT A22 A22 2155000 -6262500 METAL1
* PORT A29N A29N 2156000 -8880000 METAL1
* PORT B29 B29 2156000 -8866000 METAL1
* PORT B29N B29N 2156000 -8852000 METAL1
* PORT A29 A29 2156000 -8838000 METAL1
* PORT A25N A25N 2156000 -7464500 METAL1
* PORT B25 B25 2156000 -7450500 METAL1
* PORT B25N B25N 2156000 -7436500 METAL1
* PORT A25 A25 2156000 -7422500 METAL1
* PORT A21N A21N 2156500 -6019000 METAL1
* PORT B21 B21 2156500 -6005000 METAL1
* PORT B21N B21N 2156500 -5991000 METAL1
* PORT A21 A21 2156500 -5977000 METAL1
* PORT A28N A28N 2158000 -8608000 METAL1
* PORT B28 B28 2158000 -8594000 METAL1
* PORT B28N B28N 2158000 -8580000 METAL1
* PORT A28 A28 2158000 -8566000 METAL1
* PORT A24N A24N 2158000 -7192500 METAL1
* PORT B24 B24 2158000 -7178500 METAL1
* PORT B24N B24N 2158000 -7164500 METAL1
* PORT A24 A24 2158000 -7150500 METAL1
* PORT A20N A20N 2158500 -5747000 METAL1
* PORT B20 B20 2158500 -5733000 METAL1
* PORT B20N B20N 2158500 -5719000 METAL1
* PORT A20 A20 2158500 -5705000 METAL1
* PORT A31N A31N 2160000 -9450500 METAL1
* PORT B31 B31 2160000 -9436500 METAL1
* PORT B31N B31N 2160000 -9422500 METAL1
* PORT A31 A31 2160000 -9408500 METAL1
* PORT A27N A27N 2160000 -8035000 METAL1
* PORT B27 B27 2160000 -8021000 METAL1
* PORT B27N B27N 2160000 -8007000 METAL1
* PORT A27 A27 2160000 -7993000 METAL1
* PORT A23N A23N 2160500 -6589500 METAL1
* PORT B23 B23 2160500 -6575500 METAL1
* PORT B23N B23N 2160500 -6561500 METAL1
* PORT A23 A23 2160500 -6547500 METAL1
* PORT A14N A14N 2161000 -3437500 METAL1
* PORT B14 B14 2161000 -3423500 METAL1
* PORT B14N B14N 2161000 -3409500 METAL1
* PORT A14 A14 2161000 -3395500 METAL1
* PORT A10N A10N 2161000 -2022000 METAL1
* PORT B10 B10 2161000 -2008000 METAL1
* PORT B10N B10N 2161000 -1994000 METAL1
* PORT A10 A10 2161000 -1980000 METAL1
* PORT A18N A18N 2161500 -4899500 METAL1
* PORT B18 B18 2161500 -4885500 METAL1
* PORT B18N B18N 2161500 -4871500 METAL1
* PORT A18 A18 2161500 -4857500 METAL1
* PORT A6N A6N 2161500 -576500 METAL1
* PORT B6 B6 2161500 -562500 METAL1
* PORT B6N B6N 2161500 -548500 METAL1
* PORT A6 A6 2161500 -534500 METAL1
* PORT A13N A13N 2162500 -3152000 METAL1
* PORT B13 B13 2162500 -3138000 METAL1
* PORT B13N B13N 2162500 -3124000 METAL1
* PORT A13 A13 2162500 -3110000 METAL1
* PORT A9N A9N 2162500 -1736500 METAL1
* PORT B9 B9 2162500 -1722500 METAL1
* PORT B9N B9N 2162500 -1708500 METAL1
* PORT A9 A9 2162500 -1694500 METAL1
* PORT A17N A17N 2163000 -4614000 METAL1
* PORT B17 B17 2163000 -4600000 METAL1
* PORT B17N B17N 2163000 -4586000 METAL1
* PORT A17 A17 2163000 -4572000 METAL1
* PORT A5N A5N 2163000 -291000 METAL1
* PORT B5 B5 2163000 -277000 METAL1
* PORT B5N B5N 2163000 -263000 METAL1
* PORT A5 A5 2163000 -249000 METAL1
* PORT A12N A12N 2164500 -2880000 METAL1
* PORT B12 B12 2164500 -2866000 METAL1
* PORT B12N B12N 2164500 -2852000 METAL1
* PORT A12 A12 2164500 -2838000 METAL1
* PORT A8N A8N 2164500 -1464500 METAL1
* PORT B8 B8 2164500 -1450500 METAL1
* PORT B8N B8N 2164500 -1436500 METAL1
* PORT A8 A8 2164500 -1422500 METAL1
* PORT A16N A16N 2165000 -4342000 METAL1
* PORT B16 B16 2165000 -4328000 METAL1
* PORT B16N B16N 2165000 -4314000 METAL1
* PORT A16 A16 2165000 -4300000 METAL1
* PORT A4N A4N 2165000 -19000 METAL1
* PORT B4 B4 2165000 -5000 METAL1
* PORT B4N B4N 2165000 9000 METAL1
* PORT A4 A4 2165000 23000 METAL1
* PORT A15N A15N 2166500 -3722500 METAL1
* PORT B15 B15 2166500 -3708500 METAL1
* PORT B15N B15N 2166500 -3694500 METAL1
* PORT A15 A15 2166500 -3680500 METAL1
* PORT A11N A11N 2166500 -2307000 METAL1
* PORT B11 B11 2166500 -2293000 METAL1
* PORT B11N B11N 2166500 -2279000 METAL1
* PORT A11 A11 2166500 -2265000 METAL1
* PORT A19N A19N 2167000 -5184500 METAL1
* PORT B19 B19 2167000 -5170500 METAL1
* PORT B19N B19N 2167000 -5156500 METAL1
* PORT A19 A19 2167000 -5142500 METAL1
* PORT A7N A7N 2167000 -861500 METAL1
* PORT B7 B7 2167000 -847500 METAL1
* PORT B7N B7N 2167000 -833500 METAL1
* PORT A7 A7 2167000 -819500 METAL1
* PORT A2N A2N 2168000 828500 METAL1
* PORT B2 B2 2168000 842500 METAL1
* PORT B2N B2N 2168000 856500 METAL1
* PORT A2 A2 2168000 870500 METAL1
* PORT A1N A1N 2169500 1114000 METAL1
* PORT B1 B1 2169500 1128000 METAL1
* PORT B1N B1N 2169500 1142000 METAL1
* PORT A1 A1 2169500 1156000 METAL1
* PORT A0N A0N 2171500 1386000 METAL1
* PORT B0 B0 2171500 1400000 METAL1
* PORT B0N B0N 2171500 1414000 METAL1
* PORT A0 A0 2171500 1428000 METAL1
* PORT A3N A3N 2173500 543500 METAL1
* PORT B3 B3 2173500 557500 METAL1
* PORT B3N B3N 2173500 571500 METAL1
* PORT A3 A3 2173500 585500 METAL1
X0 VDD COUT31N 3 45 GND SUM30 SUM29 SUM28 SUM31 COUT31 A30N B30 B30N A30 A29N B29 B29N A29 A28N B28
+ B28N A28 A31N B31 B31N A31
+ four_bit_adder $T=232500 -9030500 0 0 $X=449000 $Y=-9857500
X1 VDD 3 4 46 GND SUM26 SUM25 SUM24 SUM27 45 A26N B26 B26N A26 A25N B25 B25N A25 A24N B24
+ B24N A24 A27N B27 B27N A27
+ four_bit_adder $T=232500 -7615000 0 0 $X=449000 $Y=-8442000
X2 VDD 4 5 47 GND SUM22 SUM21 SUM20 SUM23 46 A22N B22 B22N A22 A21N B21 B21N A21 A20N B20
+ B20N A20 A23N B23 B23N A23
+ four_bit_adder $T=233000 -6169500 0 0 $X=449500 $Y=-6996500
X3 VDD 8 6 48 GND SUM14 SUM13 SUM12 SUM15 50 A14N B14 B14N A14 A13N B13 B13N A13 A12N B12
+ B12N A12 A15N B15 B15N A15
+ four_bit_adder $T=239000 -3302500 0 0 $X=455500 $Y=-4129500
X4 VDD 6 7 49 GND SUM10 SUM9 SUM8 SUM11 48 A10N B10 B10N A10 A9N B9 B9N A9 A8N B8
+ B8N A8 A11N B11 B11N A11
+ four_bit_adder $T=239000 -1887000 0 0 $X=455500 $Y=-2714000
X5 VDD 5 8 50 GND SUM18 SUM17 SUM16 SUM19 47 A18N B18 B18N A18 A17N B17 B17N A17 A16N B16
+ B16N A16 A19N B19 B19N A19
+ four_bit_adder $T=239500 -4764500 0 0 $X=456000 $Y=-5591500
X6 VDD 7 9 51 GND SUM6 SUM5 SUM4 SUM7 49 A6N B6 B6N A6 A5N B5 B5N A5 A4N B4
+ B4N A4 A7N B7 B7N A7
+ four_bit_adder $T=239500 -441500 0 0 $X=456000 $Y=-1268500
X7 VDD 9 C0N C0 GND SUM2 SUM1 SUM0 SUM3 51 A2N B2 B2N A2 A1N B1 B1N A1 A0N B0
+ B0N A0 A3N B3 B3N A3
+ four_bit_adder $T=246000 963500 0 0 $X=462500 $Y=136500
.ENDS
***************************************
