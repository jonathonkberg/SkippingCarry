*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'pd433' on Mon Dec  5 2022 at 20:58:29

*
* Globals.
*
.global VDD GND

*
* MAIN CELL: Component pathname : $HOME/github/SkippingCarry/schematics/sum
*
        MN7 SUM VDD GND N$112 n L=2u W=5u
        MP7 SUM VDD VDD N$110 p L=2u W=5u
        MN6 VDD D N$101 N$107 n L=2u W=5u
        MN5 VDD B N$75 N$77 n L=2u W=5u
        MN4 N$75 A N$101 N$74 n L=2u W=5u
        MN3 VDD P N$73 N$71 n L=2u W=5u
        MN2 N$73 C__ESC1 GND N$68 n L=2u W=5u
        MP6 VDD D N$87 N$67 p L=2u W=5u
        MP5 N$88 B N$87 N$66 p L=2u W=5u
        MP4 N$87 A N$88 N$63 p L=2u W=5u
        MP3 N$88 P N$83 N$62 p L=2u W=5u
        MP2 N$83 C__ESC1 N$88 N$61 p L=2u W=5u
        MN1 N$101 C GND N$60 n L=2u W=5u
        MP1 N$88 C VDD N$59 p L=2u W=5u
*
.end
