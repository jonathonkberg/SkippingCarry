* SPICE NETLIST
***************************************

.SUBCKT i VDD IN2 IN4 IN3 IN1 OUTN OUT GND
** N=11 EP=8 IP=0 FDC=10
* PORT VDD VDD -23500 1500 METAL2
* PORT IN2 IN2 -21000 30000 METAL1
* PORT IN2 IN2 151000 58000 METAL1
* PORT IN4 IN4 -21000 44000 METAL1
* PORT IN4 IN4 151000 30000 METAL1
* PORT IN3 IN3 -21000 58000 METAL1
* PORT IN3 IN3 151000 44000 METAL1
* PORT IN1 IN1 -21000 72000 METAL1
* PORT IN1 IN1 151000 72000 METAL1
* PORT OUTN OUTN 37000 -33000 METAL1
* PORT OUT OUT 79000 -33000 METAL1
* PORT GND GND 151000 10000 METAL1
M0 GND OUTN OUT GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=90000 $Y=-12000 $D=1
M1 10 IN4 OUTN GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=113000 $Y=29000 $D=1
M2 GND IN3 10 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=43000 $D=1
M3 11 IN2 GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=57000 $D=1
M4 OUTN IN1 11 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=113000 $Y=71000 $D=1
M5 9 IN2 VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=33000 $Y=29000 $D=0
M6 OUTN IN4 9 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=43000 $D=0
M7 9 IN3 OUTN VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=57000 $D=0
M8 VDD IN1 9 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=33000 $Y=71000 $D=0
M9 VDD OUTN OUT VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=49000 $Y=-12000 $D=0
.ENDS
***************************************
.SUBCKT full_adder COUTN CN COUT C VDD SUM B A GND P AN BN
** N=21 EP=12 IP=24 FDC=44
* PORT COUTN COUTN 269500 -18000 METAL2
* PORT CN CN 286500 207500 METAL2
* PORT COUT COUT 311500 -18000 METAL1
* PORT C C 403000 190000 METAL1
* PORT VDD VDD -493000 90500 METAL1
* PORT SUM SUM -493000 29500 METAL1
* PORT B B 648000 132500 METAL1
* PORT A A 648000 160500 METAL1
* PORT GND GND 648000 98500 METAL1
* PORT P P 560000 -18000 METAL1
* PORT AN AN 648000 118500 METAL1
* PORT BN BN 648000 146500 METAL1
M0 GND 10 12 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=-121000 $Y=75000 $D=1
M1 GND 7 10 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=-118000 $Y=119000 $D=1
M2 20 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=-118000 $Y=133000 $D=1
M3 10 A 20 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=-118000 $Y=147000 $D=1
M4 GND 7 14 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=81000 $Y=76500 $D=1
M5 7 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=92000 $Y=117500 $D=1
M6 GND A 7 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=92000 $Y=131500 $D=1
M7 11 7 10 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=-177000 $Y=119000 $D=0
M8 VDD B 11 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=-177000 $Y=133000 $D=0
M9 11 A VDD VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=-177000 $Y=147000 $D=0
M10 VDD 10 12 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-162000 $Y=75000 $D=0
M11 21 B VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=31000 $Y=117500 $D=0
M12 7 A 21 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=31000 $Y=131500 $D=0
M13 VDD 7 14 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=47000 $Y=76500 $D=0
X14 VDD 12 P CN C 18 SUM GND i $T=-438000 89000 0 0 $X=-464000 $Y=54000
X15 VDD B 14 C A COUTN COUT GND i $T=232500 85000 0 0 $X=206500 $Y=50000
X16 VDD BN AN B A 19 P GND i $T=481000 88500 0 0 $X=455000 $Y=53500
.ENDS
***************************************
