* SPICE NETLIST
***************************************

.SUBCKT i VDD IN2 IN4 IN3 IN1 OUTN OUT GND
** N=11 EP=8 IP=0 FDC=10
* PORT VDD VDD -23500 1500 METAL2
* PORT IN2 IN2 -21000 30000 METAL1
* PORT IN2 IN2 151000 58000 METAL1
* PORT IN4 IN4 -21000 44000 METAL1
* PORT IN4 IN4 151000 30000 METAL1
* PORT IN3 IN3 -21000 58000 METAL1
* PORT IN3 IN3 151000 44000 METAL1
* PORT IN1 IN1 -21000 72000 METAL1
* PORT IN1 IN1 151000 72000 METAL1
* PORT OUTN OUTN 37000 -33000 METAL1
* PORT OUT OUT 79000 -33000 METAL1
* PORT GND GND 151000 10000 METAL1
M0 GND OUTN OUT GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=90000 $Y=-12000 $D=1
M1 10 IN4 OUTN GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=113000 $Y=29000 $D=1
M2 GND IN3 10 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=43000 $D=1
M3 11 IN2 GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=113000 $Y=57000 $D=1
M4 OUTN IN1 11 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=113000 $Y=71000 $D=1
M5 9 IN2 VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=33000 $Y=29000 $D=0
M6 OUTN IN4 9 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=43000 $D=0
M7 9 IN3 OUTN VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=33000 $Y=57000 $D=0
M8 VDD IN1 9 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=33000 $Y=71000 $D=0
M9 VDD OUTN OUT VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=49000 $Y=-12000 $D=0
.ENDS
***************************************
.SUBCKT full_adder COUTN CN COUT C VDD GND SUM B A P AN BN
** N=21 EP=12 IP=24 FDC=44
* PORT COUTN COUTN 269500 -18000 METAL2
* PORT CN CN 286500 207500 METAL2
* PORT COUT COUT 311500 -18000 METAL1
* PORT C C 403000 190000 METAL1
* PORT VDD VDD -493000 90500 METAL1
* PORT GND GND 648000 98500 METAL1
* PORT SUM SUM -493000 29500 METAL1
* PORT B B 648000 132500 METAL1
* PORT A A 648000 160500 METAL1
* PORT P P 560000 -18000 METAL1
* PORT AN AN 648000 118500 METAL1
* PORT BN BN 648000 146500 METAL1
M0 GND 14 16 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=-121000 $Y=75000 $D=1
M1 GND 13 14 GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=-118000 $Y=119000 $D=1
M2 20 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=-118000 $Y=133000 $D=1
M3 14 A 20 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=-118000 $Y=147000 $D=1
M4 GND 13 17 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=81000 $Y=76500 $D=1
M5 13 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=92000 $Y=117500 $D=1
M6 GND A 13 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=92000 $Y=131500 $D=1
M7 15 13 14 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=-177000 $Y=119000 $D=0
M8 VDD B 15 VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=3.1104e-12 $X=-177000 $Y=133000 $D=0
M9 15 A VDD VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=-177000 $Y=147000 $D=0
M10 VDD 14 16 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-162000 $Y=75000 $D=0
M11 21 B VDD VDD P L=1.8e-07 W=2.88e-06 AD=3.1104e-12 AS=2.3328e-12 $X=31000 $Y=117500 $D=0
M12 13 A 21 VDD P L=1.8e-07 W=2.88e-06 AD=2.3328e-12 AS=3.1104e-12 $X=31000 $Y=131500 $D=0
M13 VDD 13 17 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=47000 $Y=76500 $D=0
X14 VDD 16 P CN C 18 SUM GND i $T=-438000 89000 0 0 $X=-464000 $Y=54000
X15 VDD B 17 C A COUTN COUT GND i $T=232500 85000 0 0 $X=206500 $Y=50000
X16 VDD BN AN B A 19 P GND i $T=481000 88500 0 0 $X=455000 $Y=53500
.ENDS
***************************************
.SUBCKT four_bit_adder VDD COUTN C0N C0 GND SUM2 SUM1 SUM0 SUM3 COUT A2N B2 B2N A2 A1N B1 B1N A1 A0N B0
+ B0N A0 A3N B3 B3N A3
** N=43 EP=26 IP=56 FDC=196
* PORT VDD VDD 282000 508000 METAL2
* PORT VDD VDD 302500 -792000 METAL2
* PORT COUTN COUTN 979000 -798000 METAL2
* PORT C0N C0N 1134000 527000 METAL2
* PORT C0 C0 1250500 527000 METAL1
* PORT GND GND 1811000 519500 METAL2
* PORT GND GND 1817000 -786000 METAL2
* PORT SUM2 SUM2 218500 -224000 METAL1
* PORT SUM1 SUM1 220000 61500 METAL1
* PORT SUM0 SUM0 222000 333500 METAL1
* PORT SUM3 SUM3 224000 -509000 METAL1
* PORT COUT COUT 1021000 -798000 METAL1
* PORT A2N A2N 1894500 -135000 METAL1
* PORT B2 B2 1894500 -121000 METAL1
* PORT B2N B2N 1894500 -107000 METAL1
* PORT A2 A2 1894500 -93000 METAL1
* PORT A1N A1N 1896000 150500 METAL1
* PORT B1 B1 1896000 164500 METAL1
* PORT B1N B1N 1896000 178500 METAL1
* PORT A1 A1 1896000 192500 METAL1
* PORT A0N A0N 1898000 422500 METAL1
* PORT B0 B0 1898000 436500 METAL1
* PORT B0N B0N 1898000 450500 METAL1
* PORT A0 A0 1898000 464500 METAL1
* PORT A3N A3N 1900000 -420000 METAL1
* PORT B3 B3 1900000 -406000 METAL1
* PORT B3N B3N 1900000 -392000 METAL1
* PORT A3 A3 1900000 -378000 METAL1
M0 GND 23 24 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=1307500 $Y=-714000 $D=1
M1 41 9 GND GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=1.7496e-12 $X=1310500 $Y=-675000 $D=1
M2 42 8 41 GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12 $X=1310500 $Y=-661000 $D=1
M3 43 7 42 GND N L=1.8e-07 W=2.16e-06 AD=2.3328e-12 AS=2.3328e-12 $X=1310500 $Y=-647000 $D=1
M4 23 19 43 GND N L=1.8e-07 W=2.16e-06 AD=1.7496e-12 AS=2.3328e-12 $X=1310500 $Y=-633000 $D=1
M5 VDD 23 24 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=1266500 $Y=-714000 $D=0
M6 23 9 VDD VDD P L=1.8e-07 W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12 $X=1268500 $Y=-675000 $D=0
M7 VDD 8 23 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12 $X=1268500 $Y=-661000 $D=0
M8 23 7 VDD VDD P L=1.8e-07 W=1.44e-06 AD=1.5552e-12 AS=1.1664e-12 $X=1268500 $Y=-631000 $D=0
M9 VDD 19 23 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.5552e-12 $X=1268500 $Y=-617000 $D=0
X10 VDD 23 C0 24 18 COUTN COUT GND i $T=942000 -686000 0 0 $X=916000 $Y=-721000
X11 6 3 22 20 VDD GND SUM2 B2 A2 7 A2N B2N full_adder $T=844000 -253500 0 0 $X=349000 $Y=-273500
X12 3 4 20 21 VDD GND SUM1 B1 A1 8 A1N B1N full_adder $T=845500 32000 0 0 $X=350500 $Y=12000
X13 4 C0N 21 C0 VDD GND SUM0 B0 A0 9 A0N B0N full_adder $T=847500 304000 0 0 $X=352500 $Y=284000
X14 12 6 18 22 VDD GND SUM3 B3 A3 19 A3N B3N full_adder $T=849500 -538500 0 0 $X=354500 $Y=-558500
.ENDS
***************************************
