* File: sipo_32.pex.netlist
* Created: Thu Dec 22 00:22:57 2022
* Program "Calibre xRC"
* Version "v2012.2_36.25"
* 
.include "sipo_32.pex.netlist.pex"
.subckt SIPO_32  CLKN A3 A7 A11 A15 A19 A23 A27 A31 A0N A0 A1N A1 A2N A2 A3N A4N
+ A4 A5N A5 A6N A6 A7N A8N A8 A9N A9 A10N A10 A11N A12N A12 A13N A13 A14N A14
+ A15N A16N A16 A17N A17 A18N A18 A19N A20N A20 A21N A21 A22N A22 A23N A24N A24
+ A25N A25 A26N A26 A27N A28N A28 A29N A29 A30N A30 A31N VDD DIN GND CLK
* 
* CLK	CLK
* GND	GND
* DIN	DIN
* VDD	VDD
* A31N	A31N
* A30	A30
* A30N	A30N
* A29	A29
* A29N	A29N
* A28	A28
* A28N	A28N
* A27N	A27N
* A26	A26
* A26N	A26N
* A25	A25
* A25N	A25N
* A24	A24
* A24N	A24N
* A23N	A23N
* A22	A22
* A22N	A22N
* A21	A21
* A21N	A21N
* A20	A20
* A20N	A20N
* A19N	A19N
* A18	A18
* A18N	A18N
* A17	A17
* A17N	A17N
* A16	A16
* A16N	A16N
* A15N	A15N
* A14	A14
* A14N	A14N
* A13	A13
* A13N	A13N
* A12	A12
* A12N	A12N
* A11N	A11N
* A10	A10
* A10N	A10N
* A9	A9
* A9N	A9N
* A8	A8
* A8N	A8N
* A7N	A7N
* A6	A6
* A6N	A6N
* A5	A5
* A5N	A5N
* A4	A4
* A4N	A4N
* A3N	A3N
* A2	A2
* A2N	A2N
* A1	A1
* A1N	A1N
* A0	A0
* A0N	A0N
* A31	A31
* A27	A27
* A23	A23
* A19	A19
* A15	A15
* A11	A11
* A7	A7
* A3	A3
* CLKN	CLKN
mX0/M0 N_68_X0/M0_d N_CLKN_X0/M0_g N_X0/6_X0/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/M1 N_68_X0/M1_d N_CLKN_X0/M1_g N_X0/6_X0/M1_s N_VDD_X0/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X2/M0 N_GND_X0/X2/M0_d N_A0N_X0/X2/M0_g N_102_X0/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X2/M1 N_VDD_X0/X2/M1_d N_A0N_X0/X2/M1_g N_102_X0/X2/M1_s N_VDD_X0/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X3/M0 N_GND_X0/X3/M0_d N_A0_X0/X3/M0_g N_A0N_X0/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X3/M1 N_VDD_X0/X3/M1_d N_A0_X0/X3/M1_g N_A0N_X0/X3/M1_s N_VDD_X0/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X4/M0 N_GND_X0/X4/M0_d N_X0/5_X0/X4/M0_g N_A0_X0/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X4/M1 N_VDD_X0/X4/M1_d N_X0/5_X0/X4/M1_g N_A0_X0/X4/M1_s N_VDD_X0/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX0/X5/M0 N_GND_X0/X5/M0_d N_X0/6_X0/X5/M0_g N_X0/5_X0/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX0/X5/M1 N_VDD_X0/X5/M1_d N_X0/6_X0/X5/M1_g N_X0/5_X0/X5/M1_s N_VDD_X0/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/M0 N_69_X1/M0_d N_CLK_X1/M0_g N_X1/6_X1/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/M1 N_69_X1/M1_d N_CLK_X1/M1_g N_X1/6_X1/M1_s N_VDD_X1/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X2/M0 N_GND_X1/X2/M0_d N_A1N_X1/X2/M0_g N_68_X1/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X2/M1 N_VDD_X1/X2/M1_d N_A1N_X1/X2/M1_g N_68_X1/X2/M1_s N_VDD_X1/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X3/M0 N_GND_X1/X3/M0_d N_A1_X1/X3/M0_g N_A1N_X1/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X3/M1 N_VDD_X1/X3/M1_d N_A1_X1/X3/M1_g N_A1N_X1/X3/M1_s N_VDD_X1/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X4/M0 N_GND_X1/X4/M0_d N_X1/5_X1/X4/M0_g N_A1_X1/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X4/M1 N_VDD_X1/X4/M1_d N_X1/5_X1/X4/M1_g N_A1_X1/X4/M1_s N_VDD_X1/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX1/X5/M0 N_GND_X1/X5/M0_d N_X1/6_X1/X5/M0_g N_X1/5_X1/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX1/X5/M1 N_VDD_X1/X5/M1_d N_X1/6_X1/X5/M1_g N_X1/5_X1/X5/M1_s N_VDD_X1/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/M0 N_70_X2/M0_d N_CLKN_X2/M0_g N_X2/6_X2/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/M1 N_70_X2/M1_d N_CLKN_X2/M1_g N_X2/6_X2/M1_s N_VDD_X2/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X2/M0 N_GND_X2/X2/M0_d N_A2N_X2/X2/M0_g N_69_X2/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X2/M1 N_VDD_X2/X2/M1_d N_A2N_X2/X2/M1_g N_69_X2/X2/M1_s N_VDD_X2/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X3/M0 N_GND_X2/X3/M0_d N_A2_X2/X3/M0_g N_A2N_X2/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X3/M1 N_VDD_X2/X3/M1_d N_A2_X2/X3/M1_g N_A2N_X2/X3/M1_s N_VDD_X2/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X4/M0 N_GND_X2/X4/M0_d N_X2/5_X2/X4/M0_g N_A2_X2/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X4/M1 N_VDD_X2/X4/M1_d N_X2/5_X2/X4/M1_g N_A2_X2/X4/M1_s N_VDD_X2/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX2/X5/M0 N_GND_X2/X5/M0_d N_X2/6_X2/X5/M0_g N_X2/5_X2/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX2/X5/M1 N_VDD_X2/X5/M1_d N_X2/6_X2/X5/M1_g N_X2/5_X2/X5/M1_s N_VDD_X2/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/M0 N_71_X3/M0_d N_CLK_X3/M0_g N_X3/6_X3/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/M1 N_71_X3/M1_d N_CLK_X3/M1_g N_X3/6_X3/M1_s N_VDD_X3/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X2/M0 N_GND_X3/X2/M0_d N_A3N_X3/X2/M0_g N_70_X3/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X2/M1 N_VDD_X3/X2/M1_d N_A3N_X3/X2/M1_g N_70_X3/X2/M1_s N_VDD_X3/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X3/M0 N_GND_X3/X3/M0_d N_A3_X3/X3/M0_g N_A3N_X3/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X3/M1 N_VDD_X3/X3/M1_d N_A3_X3/X3/M1_g N_A3N_X3/X3/M1_s N_VDD_X3/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X4/M0 N_GND_X3/X4/M0_d N_X3/5_X3/X4/M0_g N_A3_X3/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X4/M1 N_VDD_X3/X4/M1_d N_X3/5_X3/X4/M1_g N_A3_X3/X4/M1_s N_VDD_X3/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX3/X5/M0 N_GND_X3/X5/M0_d N_X3/6_X3/X5/M0_g N_X3/5_X3/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX3/X5/M1 N_VDD_X3/X5/M1_d N_X3/6_X3/X5/M1_g N_X3/5_X3/X5/M1_s N_VDD_X3/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/M0 N_72_X4/M0_d N_CLKN_X4/M0_g N_X4/6_X4/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/M1 N_72_X4/M1_d N_CLKN_X4/M1_g N_X4/6_X4/M1_s N_VDD_X4/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X2/M0 N_GND_X4/X2/M0_d N_A4N_X4/X2/M0_g N_71_X4/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X2/M1 N_VDD_X4/X2/M1_d N_A4N_X4/X2/M1_g N_71_X4/X2/M1_s N_VDD_X4/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X3/M0 N_GND_X4/X3/M0_d N_A4_X4/X3/M0_g N_A4N_X4/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X3/M1 N_VDD_X4/X3/M1_d N_A4_X4/X3/M1_g N_A4N_X4/X3/M1_s N_VDD_X4/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X4/M0 N_GND_X4/X4/M0_d N_X4/5_X4/X4/M0_g N_A4_X4/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X4/M1 N_VDD_X4/X4/M1_d N_X4/5_X4/X4/M1_g N_A4_X4/X4/M1_s N_VDD_X4/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX4/X5/M0 N_GND_X4/X5/M0_d N_X4/6_X4/X5/M0_g N_X4/5_X4/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX4/X5/M1 N_VDD_X4/X5/M1_d N_X4/6_X4/X5/M1_g N_X4/5_X4/X5/M1_s N_VDD_X4/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/M0 N_73_X5/M0_d N_CLK_X5/M0_g N_X5/6_X5/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/M1 N_73_X5/M1_d N_CLK_X5/M1_g N_X5/6_X5/M1_s N_VDD_X5/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X2/M0 N_GND_X5/X2/M0_d N_A5N_X5/X2/M0_g N_72_X5/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X2/M1 N_VDD_X5/X2/M1_d N_A5N_X5/X2/M1_g N_72_X5/X2/M1_s N_VDD_X5/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X3/M0 N_GND_X5/X3/M0_d N_A5_X5/X3/M0_g N_A5N_X5/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X3/M1 N_VDD_X5/X3/M1_d N_A5_X5/X3/M1_g N_A5N_X5/X3/M1_s N_VDD_X5/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X4/M0 N_GND_X5/X4/M0_d N_X5/5_X5/X4/M0_g N_A5_X5/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X4/M1 N_VDD_X5/X4/M1_d N_X5/5_X5/X4/M1_g N_A5_X5/X4/M1_s N_VDD_X5/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX5/X5/M0 N_GND_X5/X5/M0_d N_X5/6_X5/X5/M0_g N_X5/5_X5/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX5/X5/M1 N_VDD_X5/X5/M1_d N_X5/6_X5/X5/M1_g N_X5/5_X5/X5/M1_s N_VDD_X5/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/M0 N_74_X6/M0_d N_CLKN_X6/M0_g N_X6/6_X6/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/M1 N_74_X6/M1_d N_CLKN_X6/M1_g N_X6/6_X6/M1_s N_VDD_X6/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X2/M0 N_GND_X6/X2/M0_d N_A6N_X6/X2/M0_g N_73_X6/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X2/M1 N_VDD_X6/X2/M1_d N_A6N_X6/X2/M1_g N_73_X6/X2/M1_s N_VDD_X6/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X3/M0 N_GND_X6/X3/M0_d N_A6_X6/X3/M0_g N_A6N_X6/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X3/M1 N_VDD_X6/X3/M1_d N_A6_X6/X3/M1_g N_A6N_X6/X3/M1_s N_VDD_X6/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X4/M0 N_GND_X6/X4/M0_d N_X6/5_X6/X4/M0_g N_A6_X6/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X4/M1 N_VDD_X6/X4/M1_d N_X6/5_X6/X4/M1_g N_A6_X6/X4/M1_s N_VDD_X6/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX6/X5/M0 N_GND_X6/X5/M0_d N_X6/6_X6/X5/M0_g N_X6/5_X6/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX6/X5/M1 N_VDD_X6/X5/M1_d N_X6/6_X6/X5/M1_g N_X6/5_X6/X5/M1_s N_VDD_X6/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/M0 N_75_X7/M0_d N_CLK_X7/M0_g N_X7/6_X7/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/M1 N_75_X7/M1_d N_CLK_X7/M1_g N_X7/6_X7/M1_s N_VDD_X7/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X2/M0 N_GND_X7/X2/M0_d N_A7N_X7/X2/M0_g N_74_X7/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X2/M1 N_VDD_X7/X2/M1_d N_A7N_X7/X2/M1_g N_74_X7/X2/M1_s N_VDD_X7/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X3/M0 N_GND_X7/X3/M0_d N_A7_X7/X3/M0_g N_A7N_X7/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X3/M1 N_VDD_X7/X3/M1_d N_A7_X7/X3/M1_g N_A7N_X7/X3/M1_s N_VDD_X7/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X4/M0 N_GND_X7/X4/M0_d N_X7/5_X7/X4/M0_g N_A7_X7/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X4/M1 N_VDD_X7/X4/M1_d N_X7/5_X7/X4/M1_g N_A7_X7/X4/M1_s N_VDD_X7/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX7/X5/M0 N_GND_X7/X5/M0_d N_X7/6_X7/X5/M0_g N_X7/5_X7/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX7/X5/M1 N_VDD_X7/X5/M1_d N_X7/6_X7/X5/M1_g N_X7/5_X7/X5/M1_s N_VDD_X7/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX8/M0 N_76_X8/M0_d N_CLKN_X8/M0_g N_X8/6_X8/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX8/M1 N_76_X8/M1_d N_CLKN_X8/M1_g N_X8/6_X8/M1_s N_VDD_X8/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX8/X2/M0 N_GND_X8/X2/M0_d N_A8N_X8/X2/M0_g N_75_X8/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX8/X2/M1 N_VDD_X8/X2/M1_d N_A8N_X8/X2/M1_g N_75_X8/X2/M1_s N_VDD_X8/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX8/X3/M0 N_GND_X8/X3/M0_d N_A8_X8/X3/M0_g N_A8N_X8/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX8/X3/M1 N_VDD_X8/X3/M1_d N_A8_X8/X3/M1_g N_A8N_X8/X3/M1_s N_VDD_X8/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX8/X4/M0 N_GND_X8/X4/M0_d N_X8/5_X8/X4/M0_g N_A8_X8/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX8/X4/M1 N_VDD_X8/X4/M1_d N_X8/5_X8/X4/M1_g N_A8_X8/X4/M1_s N_VDD_X8/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX8/X5/M0 N_GND_X8/X5/M0_d N_X8/6_X8/X5/M0_g N_X8/5_X8/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX8/X5/M1 N_VDD_X8/X5/M1_d N_X8/6_X8/X5/M1_g N_X8/5_X8/X5/M1_s N_VDD_X8/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX9/M0 N_77_X9/M0_d N_CLK_X9/M0_g N_X9/6_X9/M0_s N_GND_X0/X2/M0_b n L=1.8e-07
+ W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX9/M1 N_77_X9/M1_d N_CLK_X9/M1_g N_X9/6_X9/M1_s N_VDD_X9/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX9/X2/M0 N_GND_X9/X2/M0_d N_A9N_X9/X2/M0_g N_76_X9/X2/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX9/X2/M1 N_VDD_X9/X2/M1_d N_A9N_X9/X2/M1_g N_76_X9/X2/M1_s N_VDD_X9/X2/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX9/X3/M0 N_GND_X9/X3/M0_d N_A9_X9/X3/M0_g N_A9N_X9/X3/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX9/X3/M1 N_VDD_X9/X3/M1_d N_A9_X9/X3/M1_g N_A9N_X9/X3/M1_s N_VDD_X9/X3/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX9/X4/M0 N_GND_X9/X4/M0_d N_X9/5_X9/X4/M0_g N_A9_X9/X4/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX9/X4/M1 N_VDD_X9/X4/M1_d N_X9/5_X9/X4/M1_g N_A9_X9/X4/M1_s N_VDD_X9/X4/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX9/X5/M0 N_GND_X9/X5/M0_d N_X9/6_X9/X5/M0_g N_X9/5_X9/X5/M0_s N_GND_X0/X2/M0_b
+ n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX9/X5/M1 N_VDD_X9/X5/M1_d N_X9/6_X9/X5/M1_g N_X9/5_X9/X5/M1_s N_VDD_X9/X5/M1_b
+ p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX10/M0 N_78_X10/M0_d N_CLKN_X10/M0_g N_X10/6_X10/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX10/M1 N_78_X10/M1_d N_CLKN_X10/M1_g N_X10/6_X10/M1_s N_VDD_X10/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX10/X2/M0 N_GND_X10/X2/M0_d N_A10N_X10/X2/M0_g N_77_X10/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX10/X2/M1 N_VDD_X10/X2/M1_d N_A10N_X10/X2/M1_g N_77_X10/X2/M1_s
+ N_VDD_X10/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX10/X3/M0 N_GND_X10/X3/M0_d N_A10_X10/X3/M0_g N_A10N_X10/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX10/X3/M1 N_VDD_X10/X3/M1_d N_A10_X10/X3/M1_g N_A10N_X10/X3/M1_s
+ N_VDD_X10/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX10/X4/M0 N_GND_X10/X4/M0_d N_X10/5_X10/X4/M0_g N_A10_X10/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX10/X4/M1 N_VDD_X10/X4/M1_d N_X10/5_X10/X4/M1_g N_A10_X10/X4/M1_s
+ N_VDD_X10/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX10/X5/M0 N_GND_X10/X5/M0_d N_X10/6_X10/X5/M0_g N_X10/5_X10/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX10/X5/M1 N_VDD_X10/X5/M1_d N_X10/6_X10/X5/M1_g N_X10/5_X10/X5/M1_s
+ N_VDD_X10/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX11/M0 N_79_X11/M0_d N_CLK_X11/M0_g N_X11/6_X11/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX11/M1 N_79_X11/M1_d N_CLK_X11/M1_g N_X11/6_X11/M1_s N_VDD_X11/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX11/X2/M0 N_GND_X11/X2/M0_d N_A11N_X11/X2/M0_g N_78_X11/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX11/X2/M1 N_VDD_X11/X2/M1_d N_A11N_X11/X2/M1_g N_78_X11/X2/M1_s
+ N_VDD_X11/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX11/X3/M0 N_GND_X11/X3/M0_d N_A11_X11/X3/M0_g N_A11N_X11/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX11/X3/M1 N_VDD_X11/X3/M1_d N_A11_X11/X3/M1_g N_A11N_X11/X3/M1_s
+ N_VDD_X11/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX11/X4/M0 N_GND_X11/X4/M0_d N_X11/5_X11/X4/M0_g N_A11_X11/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX11/X4/M1 N_VDD_X11/X4/M1_d N_X11/5_X11/X4/M1_g N_A11_X11/X4/M1_s
+ N_VDD_X11/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX11/X5/M0 N_GND_X11/X5/M0_d N_X11/6_X11/X5/M0_g N_X11/5_X11/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX11/X5/M1 N_VDD_X11/X5/M1_d N_X11/6_X11/X5/M1_g N_X11/5_X11/X5/M1_s
+ N_VDD_X11/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX12/M0 N_80_X12/M0_d N_CLKN_X12/M0_g N_X12/6_X12/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX12/M1 N_80_X12/M1_d N_CLKN_X12/M1_g N_X12/6_X12/M1_s N_VDD_X12/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX12/X2/M0 N_GND_X12/X2/M0_d N_A12N_X12/X2/M0_g N_79_X12/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX12/X2/M1 N_VDD_X12/X2/M1_d N_A12N_X12/X2/M1_g N_79_X12/X2/M1_s
+ N_VDD_X12/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX12/X3/M0 N_GND_X12/X3/M0_d N_A12_X12/X3/M0_g N_A12N_X12/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX12/X3/M1 N_VDD_X12/X3/M1_d N_A12_X12/X3/M1_g N_A12N_X12/X3/M1_s
+ N_VDD_X12/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX12/X4/M0 N_GND_X12/X4/M0_d N_X12/5_X12/X4/M0_g N_A12_X12/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX12/X4/M1 N_VDD_X12/X4/M1_d N_X12/5_X12/X4/M1_g N_A12_X12/X4/M1_s
+ N_VDD_X12/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX12/X5/M0 N_GND_X12/X5/M0_d N_X12/6_X12/X5/M0_g N_X12/5_X12/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX12/X5/M1 N_VDD_X12/X5/M1_d N_X12/6_X12/X5/M1_g N_X12/5_X12/X5/M1_s
+ N_VDD_X12/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX13/M0 N_81_X13/M0_d N_CLK_X13/M0_g N_X13/6_X13/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX13/M1 N_81_X13/M1_d N_CLK_X13/M1_g N_X13/6_X13/M1_s N_VDD_X13/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX13/X2/M0 N_GND_X13/X2/M0_d N_A13N_X13/X2/M0_g N_80_X13/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX13/X2/M1 N_VDD_X13/X2/M1_d N_A13N_X13/X2/M1_g N_80_X13/X2/M1_s
+ N_VDD_X13/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX13/X3/M0 N_GND_X13/X3/M0_d N_A13_X13/X3/M0_g N_A13N_X13/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX13/X3/M1 N_VDD_X13/X3/M1_d N_A13_X13/X3/M1_g N_A13N_X13/X3/M1_s
+ N_VDD_X13/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX13/X4/M0 N_GND_X13/X4/M0_d N_X13/5_X13/X4/M0_g N_A13_X13/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX13/X4/M1 N_VDD_X13/X4/M1_d N_X13/5_X13/X4/M1_g N_A13_X13/X4/M1_s
+ N_VDD_X13/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX13/X5/M0 N_GND_X13/X5/M0_d N_X13/6_X13/X5/M0_g N_X13/5_X13/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX13/X5/M1 N_VDD_X13/X5/M1_d N_X13/6_X13/X5/M1_g N_X13/5_X13/X5/M1_s
+ N_VDD_X13/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX14/M0 N_82_X14/M0_d N_CLKN_X14/M0_g N_X14/6_X14/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX14/M1 N_82_X14/M1_d N_CLKN_X14/M1_g N_X14/6_X14/M1_s N_VDD_X14/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX14/X2/M0 N_GND_X14/X2/M0_d N_A14N_X14/X2/M0_g N_81_X14/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX14/X2/M1 N_VDD_X14/X2/M1_d N_A14N_X14/X2/M1_g N_81_X14/X2/M1_s
+ N_VDD_X14/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX14/X3/M0 N_GND_X14/X3/M0_d N_A14_X14/X3/M0_g N_A14N_X14/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX14/X3/M1 N_VDD_X14/X3/M1_d N_A14_X14/X3/M1_g N_A14N_X14/X3/M1_s
+ N_VDD_X14/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX14/X4/M0 N_GND_X14/X4/M0_d N_X14/5_X14/X4/M0_g N_A14_X14/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX14/X4/M1 N_VDD_X14/X4/M1_d N_X14/5_X14/X4/M1_g N_A14_X14/X4/M1_s
+ N_VDD_X14/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX14/X5/M0 N_GND_X14/X5/M0_d N_X14/6_X14/X5/M0_g N_X14/5_X14/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX14/X5/M1 N_VDD_X14/X5/M1_d N_X14/6_X14/X5/M1_g N_X14/5_X14/X5/M1_s
+ N_VDD_X14/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX15/M0 N_83_X15/M0_d N_CLK_X15/M0_g N_X15/6_X15/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX15/M1 N_83_X15/M1_d N_CLK_X15/M1_g N_X15/6_X15/M1_s N_VDD_X15/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX15/X2/M0 N_GND_X15/X2/M0_d N_A15N_X15/X2/M0_g N_82_X15/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX15/X2/M1 N_VDD_X15/X2/M1_d N_A15N_X15/X2/M1_g N_82_X15/X2/M1_s
+ N_VDD_X15/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX15/X3/M0 N_GND_X15/X3/M0_d N_A15_X15/X3/M0_g N_A15N_X15/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX15/X3/M1 N_VDD_X15/X3/M1_d N_A15_X15/X3/M1_g N_A15N_X15/X3/M1_s
+ N_VDD_X15/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX15/X4/M0 N_GND_X15/X4/M0_d N_X15/5_X15/X4/M0_g N_A15_X15/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX15/X4/M1 N_VDD_X15/X4/M1_d N_X15/5_X15/X4/M1_g N_A15_X15/X4/M1_s
+ N_VDD_X15/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX15/X5/M0 N_GND_X15/X5/M0_d N_X15/6_X15/X5/M0_g N_X15/5_X15/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX15/X5/M1 N_VDD_X15/X5/M1_d N_X15/6_X15/X5/M1_g N_X15/5_X15/X5/M1_s
+ N_VDD_X15/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX16/M0 N_84_X16/M0_d N_CLKN_X16/M0_g N_X16/6_X16/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX16/M1 N_84_X16/M1_d N_CLKN_X16/M1_g N_X16/6_X16/M1_s N_VDD_X16/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX16/X2/M0 N_GND_X16/X2/M0_d N_A16N_X16/X2/M0_g N_83_X16/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX16/X2/M1 N_VDD_X16/X2/M1_d N_A16N_X16/X2/M1_g N_83_X16/X2/M1_s
+ N_VDD_X16/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX16/X3/M0 N_GND_X16/X3/M0_d N_A16_X16/X3/M0_g N_A16N_X16/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX16/X3/M1 N_VDD_X16/X3/M1_d N_A16_X16/X3/M1_g N_A16N_X16/X3/M1_s
+ N_VDD_X16/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX16/X4/M0 N_GND_X16/X4/M0_d N_X16/5_X16/X4/M0_g N_A16_X16/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX16/X4/M1 N_VDD_X16/X4/M1_d N_X16/5_X16/X4/M1_g N_A16_X16/X4/M1_s
+ N_VDD_X16/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX16/X5/M0 N_GND_X16/X5/M0_d N_X16/6_X16/X5/M0_g N_X16/5_X16/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX16/X5/M1 N_VDD_X16/X5/M1_d N_X16/6_X16/X5/M1_g N_X16/5_X16/X5/M1_s
+ N_VDD_X16/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX17/M0 N_85_X17/M0_d N_CLK_X17/M0_g N_X17/6_X17/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX17/M1 N_85_X17/M1_d N_CLK_X17/M1_g N_X17/6_X17/M1_s N_VDD_X17/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX17/X2/M0 N_GND_X17/X2/M0_d N_A17N_X17/X2/M0_g N_84_X17/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX17/X2/M1 N_VDD_X17/X2/M1_d N_A17N_X17/X2/M1_g N_84_X17/X2/M1_s
+ N_VDD_X17/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX17/X3/M0 N_GND_X17/X3/M0_d N_A17_X17/X3/M0_g N_A17N_X17/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX17/X3/M1 N_VDD_X17/X3/M1_d N_A17_X17/X3/M1_g N_A17N_X17/X3/M1_s
+ N_VDD_X17/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX17/X4/M0 N_GND_X17/X4/M0_d N_X17/5_X17/X4/M0_g N_A17_X17/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX17/X4/M1 N_VDD_X17/X4/M1_d N_X17/5_X17/X4/M1_g N_A17_X17/X4/M1_s
+ N_VDD_X17/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX17/X5/M0 N_GND_X17/X5/M0_d N_X17/6_X17/X5/M0_g N_X17/5_X17/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX17/X5/M1 N_VDD_X17/X5/M1_d N_X17/6_X17/X5/M1_g N_X17/5_X17/X5/M1_s
+ N_VDD_X17/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX18/M0 N_86_X18/M0_d N_CLKN_X18/M0_g N_X18/6_X18/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX18/M1 N_86_X18/M1_d N_CLKN_X18/M1_g N_X18/6_X18/M1_s N_VDD_X18/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX18/X2/M0 N_GND_X18/X2/M0_d N_A18N_X18/X2/M0_g N_85_X18/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX18/X2/M1 N_VDD_X18/X2/M1_d N_A18N_X18/X2/M1_g N_85_X18/X2/M1_s
+ N_VDD_X18/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX18/X3/M0 N_GND_X18/X3/M0_d N_A18_X18/X3/M0_g N_A18N_X18/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX18/X3/M1 N_VDD_X18/X3/M1_d N_A18_X18/X3/M1_g N_A18N_X18/X3/M1_s
+ N_VDD_X18/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX18/X4/M0 N_GND_X18/X4/M0_d N_X18/5_X18/X4/M0_g N_A18_X18/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX18/X4/M1 N_VDD_X18/X4/M1_d N_X18/5_X18/X4/M1_g N_A18_X18/X4/M1_s
+ N_VDD_X18/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX18/X5/M0 N_GND_X18/X5/M0_d N_X18/6_X18/X5/M0_g N_X18/5_X18/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX18/X5/M1 N_VDD_X18/X5/M1_d N_X18/6_X18/X5/M1_g N_X18/5_X18/X5/M1_s
+ N_VDD_X18/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX19/M0 N_87_X19/M0_d N_CLK_X19/M0_g N_X19/6_X19/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX19/M1 N_87_X19/M1_d N_CLK_X19/M1_g N_X19/6_X19/M1_s N_VDD_X19/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX19/X2/M0 N_GND_X19/X2/M0_d N_A19N_X19/X2/M0_g N_86_X19/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX19/X2/M1 N_VDD_X19/X2/M1_d N_A19N_X19/X2/M1_g N_86_X19/X2/M1_s
+ N_VDD_X19/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX19/X3/M0 N_GND_X19/X3/M0_d N_A19_X19/X3/M0_g N_A19N_X19/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX19/X3/M1 N_VDD_X19/X3/M1_d N_A19_X19/X3/M1_g N_A19N_X19/X3/M1_s
+ N_VDD_X19/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX19/X4/M0 N_GND_X19/X4/M0_d N_X19/5_X19/X4/M0_g N_A19_X19/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX19/X4/M1 N_VDD_X19/X4/M1_d N_X19/5_X19/X4/M1_g N_A19_X19/X4/M1_s
+ N_VDD_X19/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX19/X5/M0 N_GND_X19/X5/M0_d N_X19/6_X19/X5/M0_g N_X19/5_X19/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX19/X5/M1 N_VDD_X19/X5/M1_d N_X19/6_X19/X5/M1_g N_X19/5_X19/X5/M1_s
+ N_VDD_X19/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX20/M0 N_88_X20/M0_d N_CLKN_X20/M0_g N_X20/6_X20/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX20/M1 N_88_X20/M1_d N_CLKN_X20/M1_g N_X20/6_X20/M1_s N_VDD_X20/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX20/X2/M0 N_GND_X20/X2/M0_d N_A20N_X20/X2/M0_g N_87_X20/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX20/X2/M1 N_VDD_X20/X2/M1_d N_A20N_X20/X2/M1_g N_87_X20/X2/M1_s
+ N_VDD_X20/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX20/X3/M0 N_GND_X20/X3/M0_d N_A20_X20/X3/M0_g N_A20N_X20/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX20/X3/M1 N_VDD_X20/X3/M1_d N_A20_X20/X3/M1_g N_A20N_X20/X3/M1_s
+ N_VDD_X20/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX20/X4/M0 N_GND_X20/X4/M0_d N_X20/5_X20/X4/M0_g N_A20_X20/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX20/X4/M1 N_VDD_X20/X4/M1_d N_X20/5_X20/X4/M1_g N_A20_X20/X4/M1_s
+ N_VDD_X20/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX20/X5/M0 N_GND_X20/X5/M0_d N_X20/6_X20/X5/M0_g N_X20/5_X20/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX20/X5/M1 N_VDD_X20/X5/M1_d N_X20/6_X20/X5/M1_g N_X20/5_X20/X5/M1_s
+ N_VDD_X20/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX21/M0 N_89_X21/M0_d N_CLK_X21/M0_g N_X21/6_X21/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX21/M1 N_89_X21/M1_d N_CLK_X21/M1_g N_X21/6_X21/M1_s N_VDD_X21/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX21/X2/M0 N_GND_X21/X2/M0_d N_A21N_X21/X2/M0_g N_88_X21/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX21/X2/M1 N_VDD_X21/X2/M1_d N_A21N_X21/X2/M1_g N_88_X21/X2/M1_s
+ N_VDD_X21/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX21/X3/M0 N_GND_X21/X3/M0_d N_A21_X21/X3/M0_g N_A21N_X21/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX21/X3/M1 N_VDD_X21/X3/M1_d N_A21_X21/X3/M1_g N_A21N_X21/X3/M1_s
+ N_VDD_X21/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX21/X4/M0 N_GND_X21/X4/M0_d N_X21/5_X21/X4/M0_g N_A21_X21/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX21/X4/M1 N_VDD_X21/X4/M1_d N_X21/5_X21/X4/M1_g N_A21_X21/X4/M1_s
+ N_VDD_X21/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX21/X5/M0 N_GND_X21/X5/M0_d N_X21/6_X21/X5/M0_g N_X21/5_X21/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX21/X5/M1 N_VDD_X21/X5/M1_d N_X21/6_X21/X5/M1_g N_X21/5_X21/X5/M1_s
+ N_VDD_X21/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX22/M0 N_90_X22/M0_d N_CLKN_X22/M0_g N_X22/6_X22/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX22/M1 N_90_X22/M1_d N_CLKN_X22/M1_g N_X22/6_X22/M1_s N_VDD_X22/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX22/X2/M0 N_GND_X22/X2/M0_d N_A22N_X22/X2/M0_g N_89_X22/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX22/X2/M1 N_VDD_X22/X2/M1_d N_A22N_X22/X2/M1_g N_89_X22/X2/M1_s
+ N_VDD_X22/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX22/X3/M0 N_GND_X22/X3/M0_d N_A22_X22/X3/M0_g N_A22N_X22/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX22/X3/M1 N_VDD_X22/X3/M1_d N_A22_X22/X3/M1_g N_A22N_X22/X3/M1_s
+ N_VDD_X22/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX22/X4/M0 N_GND_X22/X4/M0_d N_X22/5_X22/X4/M0_g N_A22_X22/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX22/X4/M1 N_VDD_X22/X4/M1_d N_X22/5_X22/X4/M1_g N_A22_X22/X4/M1_s
+ N_VDD_X22/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX22/X5/M0 N_GND_X22/X5/M0_d N_X22/6_X22/X5/M0_g N_X22/5_X22/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX22/X5/M1 N_VDD_X22/X5/M1_d N_X22/6_X22/X5/M1_g N_X22/5_X22/X5/M1_s
+ N_VDD_X22/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX23/M0 N_91_X23/M0_d N_CLK_X23/M0_g N_X23/6_X23/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX23/M1 N_91_X23/M1_d N_CLK_X23/M1_g N_X23/6_X23/M1_s N_VDD_X23/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX23/X2/M0 N_GND_X23/X2/M0_d N_A23N_X23/X2/M0_g N_90_X23/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX23/X2/M1 N_VDD_X23/X2/M1_d N_A23N_X23/X2/M1_g N_90_X23/X2/M1_s
+ N_VDD_X23/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX23/X3/M0 N_GND_X23/X3/M0_d N_A23_X23/X3/M0_g N_A23N_X23/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX23/X3/M1 N_VDD_X23/X3/M1_d N_A23_X23/X3/M1_g N_A23N_X23/X3/M1_s
+ N_VDD_X23/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX23/X4/M0 N_GND_X23/X4/M0_d N_X23/5_X23/X4/M0_g N_A23_X23/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX23/X4/M1 N_VDD_X23/X4/M1_d N_X23/5_X23/X4/M1_g N_A23_X23/X4/M1_s
+ N_VDD_X23/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX23/X5/M0 N_GND_X23/X5/M0_d N_X23/6_X23/X5/M0_g N_X23/5_X23/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX23/X5/M1 N_VDD_X23/X5/M1_d N_X23/6_X23/X5/M1_g N_X23/5_X23/X5/M1_s
+ N_VDD_X23/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX24/M0 N_92_X24/M0_d N_CLKN_X24/M0_g N_X24/6_X24/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX24/M1 N_92_X24/M1_d N_CLKN_X24/M1_g N_X24/6_X24/M1_s N_VDD_X24/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX24/X2/M0 N_GND_X24/X2/M0_d N_A24N_X24/X2/M0_g N_91_X24/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX24/X2/M1 N_VDD_X24/X2/M1_d N_A24N_X24/X2/M1_g N_91_X24/X2/M1_s
+ N_VDD_X24/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX24/X3/M0 N_GND_X24/X3/M0_d N_A24_X24/X3/M0_g N_A24N_X24/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX24/X3/M1 N_VDD_X24/X3/M1_d N_A24_X24/X3/M1_g N_A24N_X24/X3/M1_s
+ N_VDD_X24/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX24/X4/M0 N_GND_X24/X4/M0_d N_X24/5_X24/X4/M0_g N_A24_X24/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX24/X4/M1 N_VDD_X24/X4/M1_d N_X24/5_X24/X4/M1_g N_A24_X24/X4/M1_s
+ N_VDD_X24/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX24/X5/M0 N_GND_X24/X5/M0_d N_X24/6_X24/X5/M0_g N_X24/5_X24/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX24/X5/M1 N_VDD_X24/X5/M1_d N_X24/6_X24/X5/M1_g N_X24/5_X24/X5/M1_s
+ N_VDD_X24/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX25/M0 N_93_X25/M0_d N_CLK_X25/M0_g N_X25/6_X25/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX25/M1 N_93_X25/M1_d N_CLK_X25/M1_g N_X25/6_X25/M1_s N_VDD_X25/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX25/X2/M0 N_GND_X25/X2/M0_d N_A25N_X25/X2/M0_g N_92_X25/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX25/X2/M1 N_VDD_X25/X2/M1_d N_A25N_X25/X2/M1_g N_92_X25/X2/M1_s
+ N_VDD_X25/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX25/X3/M0 N_GND_X25/X3/M0_d N_A25_X25/X3/M0_g N_A25N_X25/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX25/X3/M1 N_VDD_X25/X3/M1_d N_A25_X25/X3/M1_g N_A25N_X25/X3/M1_s
+ N_VDD_X25/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX25/X4/M0 N_GND_X25/X4/M0_d N_X25/5_X25/X4/M0_g N_A25_X25/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX25/X4/M1 N_VDD_X25/X4/M1_d N_X25/5_X25/X4/M1_g N_A25_X25/X4/M1_s
+ N_VDD_X25/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX25/X5/M0 N_GND_X25/X5/M0_d N_X25/6_X25/X5/M0_g N_X25/5_X25/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX25/X5/M1 N_VDD_X25/X5/M1_d N_X25/6_X25/X5/M1_g N_X25/5_X25/X5/M1_s
+ N_VDD_X25/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX26/M0 N_94_X26/M0_d N_CLKN_X26/M0_g N_X26/6_X26/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX26/M1 N_94_X26/M1_d N_CLKN_X26/M1_g N_X26/6_X26/M1_s N_VDD_X26/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX26/X2/M0 N_GND_X26/X2/M0_d N_A26N_X26/X2/M0_g N_93_X26/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX26/X2/M1 N_VDD_X26/X2/M1_d N_A26N_X26/X2/M1_g N_93_X26/X2/M1_s
+ N_VDD_X26/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX26/X3/M0 N_GND_X26/X3/M0_d N_A26_X26/X3/M0_g N_A26N_X26/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX26/X3/M1 N_VDD_X26/X3/M1_d N_A26_X26/X3/M1_g N_A26N_X26/X3/M1_s
+ N_VDD_X26/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX26/X4/M0 N_GND_X26/X4/M0_d N_X26/5_X26/X4/M0_g N_A26_X26/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX26/X4/M1 N_VDD_X26/X4/M1_d N_X26/5_X26/X4/M1_g N_A26_X26/X4/M1_s
+ N_VDD_X26/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX26/X5/M0 N_GND_X26/X5/M0_d N_X26/6_X26/X5/M0_g N_X26/5_X26/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX26/X5/M1 N_VDD_X26/X5/M1_d N_X26/6_X26/X5/M1_g N_X26/5_X26/X5/M1_s
+ N_VDD_X26/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX27/M0 N_95_X27/M0_d N_CLK_X27/M0_g N_X27/6_X27/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX27/M1 N_95_X27/M1_d N_CLK_X27/M1_g N_X27/6_X27/M1_s N_VDD_X27/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX27/X2/M0 N_GND_X27/X2/M0_d N_A27N_X27/X2/M0_g N_94_X27/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX27/X2/M1 N_VDD_X27/X2/M1_d N_A27N_X27/X2/M1_g N_94_X27/X2/M1_s
+ N_VDD_X27/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX27/X3/M0 N_GND_X27/X3/M0_d N_A27_X27/X3/M0_g N_A27N_X27/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX27/X3/M1 N_VDD_X27/X3/M1_d N_A27_X27/X3/M1_g N_A27N_X27/X3/M1_s
+ N_VDD_X27/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX27/X4/M0 N_GND_X27/X4/M0_d N_X27/5_X27/X4/M0_g N_A27_X27/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX27/X4/M1 N_VDD_X27/X4/M1_d N_X27/5_X27/X4/M1_g N_A27_X27/X4/M1_s
+ N_VDD_X27/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX27/X5/M0 N_GND_X27/X5/M0_d N_X27/6_X27/X5/M0_g N_X27/5_X27/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX27/X5/M1 N_VDD_X27/X5/M1_d N_X27/6_X27/X5/M1_g N_X27/5_X27/X5/M1_s
+ N_VDD_X27/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX28/M0 N_96_X28/M0_d N_CLKN_X28/M0_g N_X28/6_X28/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX28/M1 N_96_X28/M1_d N_CLKN_X28/M1_g N_X28/6_X28/M1_s N_VDD_X28/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX28/X2/M0 N_GND_X28/X2/M0_d N_A28N_X28/X2/M0_g N_95_X28/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX28/X2/M1 N_VDD_X28/X2/M1_d N_A28N_X28/X2/M1_g N_95_X28/X2/M1_s
+ N_VDD_X28/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX28/X3/M0 N_GND_X28/X3/M0_d N_A28_X28/X3/M0_g N_A28N_X28/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX28/X3/M1 N_VDD_X28/X3/M1_d N_A28_X28/X3/M1_g N_A28N_X28/X3/M1_s
+ N_VDD_X28/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX28/X4/M0 N_GND_X28/X4/M0_d N_X28/5_X28/X4/M0_g N_A28_X28/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX28/X4/M1 N_VDD_X28/X4/M1_d N_X28/5_X28/X4/M1_g N_A28_X28/X4/M1_s
+ N_VDD_X28/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX28/X5/M0 N_GND_X28/X5/M0_d N_X28/6_X28/X5/M0_g N_X28/5_X28/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX28/X5/M1 N_VDD_X28/X5/M1_d N_X28/6_X28/X5/M1_g N_X28/5_X28/X5/M1_s
+ N_VDD_X28/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX29/M0 N_97_X29/M0_d N_CLK_X29/M0_g N_X29/6_X29/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX29/M1 N_97_X29/M1_d N_CLK_X29/M1_g N_X29/6_X29/M1_s N_VDD_X29/M1_b p L=1.8e-07
+ W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX29/X2/M0 N_GND_X29/X2/M0_d N_A29N_X29/X2/M0_g N_96_X29/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX29/X2/M1 N_VDD_X29/X2/M1_d N_A29N_X29/X2/M1_g N_96_X29/X2/M1_s
+ N_VDD_X29/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX29/X3/M0 N_GND_X29/X3/M0_d N_A29_X29/X3/M0_g N_A29N_X29/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX29/X3/M1 N_VDD_X29/X3/M1_d N_A29_X29/X3/M1_g N_A29N_X29/X3/M1_s
+ N_VDD_X29/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX29/X4/M0 N_GND_X29/X4/M0_d N_X29/5_X29/X4/M0_g N_A29_X29/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX29/X4/M1 N_VDD_X29/X4/M1_d N_X29/5_X29/X4/M1_g N_A29_X29/X4/M1_s
+ N_VDD_X29/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX29/X5/M0 N_GND_X29/X5/M0_d N_X29/6_X29/X5/M0_g N_X29/5_X29/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX29/X5/M1 N_VDD_X29/X5/M1_d N_X29/6_X29/X5/M1_g N_X29/5_X29/X5/M1_s
+ N_VDD_X29/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX30/M0 N_98_X30/M0_d N_CLKN_X30/M0_g N_X30/6_X30/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX30/M1 N_98_X30/M1_d N_CLKN_X30/M1_g N_X30/6_X30/M1_s N_VDD_X30/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX30/X2/M0 N_GND_X30/X2/M0_d N_A30N_X30/X2/M0_g N_97_X30/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX30/X2/M1 N_VDD_X30/X2/M1_d N_A30N_X30/X2/M1_g N_97_X30/X2/M1_s
+ N_VDD_X30/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX30/X3/M0 N_GND_X30/X3/M0_d N_A30_X30/X3/M0_g N_A30N_X30/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX30/X3/M1 N_VDD_X30/X3/M1_d N_A30_X30/X3/M1_g N_A30N_X30/X3/M1_s
+ N_VDD_X30/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX30/X4/M0 N_GND_X30/X4/M0_d N_X30/5_X30/X4/M0_g N_A30_X30/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX30/X4/M1 N_VDD_X30/X4/M1_d N_X30/5_X30/X4/M1_g N_A30_X30/X4/M1_s
+ N_VDD_X30/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX30/X5/M0 N_GND_X30/X5/M0_d N_X30/6_X30/X5/M0_g N_X30/5_X30/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX30/X5/M1 N_VDD_X30/X5/M1_d N_X30/6_X30/X5/M1_g N_X30/5_X30/X5/M1_s
+ N_VDD_X30/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX31/M0 N_DIN_X31/M0_d N_CLK_X31/M0_g N_X31/6_X31/M0_s N_GND_X0/X2/M0_b n
+ L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX31/M1 N_DIN_X31/M1_d N_CLK_X31/M1_g N_X31/6_X31/M1_s N_VDD_X31/M1_b p
+ L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX31/X2/M0 N_GND_X31/X2/M0_d N_A31N_X31/X2/M0_g N_98_X31/X2/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX31/X2/M1 N_VDD_X31/X2/M1_d N_A31N_X31/X2/M1_g N_98_X31/X2/M1_s
+ N_VDD_X31/X2/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX31/X3/M0 N_GND_X31/X3/M0_d N_A31_X31/X3/M0_g N_A31N_X31/X3/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX31/X3/M1 N_VDD_X31/X3/M1_d N_A31_X31/X3/M1_g N_A31N_X31/X3/M1_s
+ N_VDD_X31/X3/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX31/X4/M0 N_GND_X31/X4/M0_d N_X31/5_X31/X4/M0_g N_A31_X31/X4/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX31/X4/M1 N_VDD_X31/X4/M1_d N_X31/5_X31/X4/M1_g N_A31_X31/X4/M1_s
+ N_VDD_X31/X4/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
mX31/X5/M0 N_GND_X31/X5/M0_d N_X31/6_X31/X5/M0_g N_X31/5_X31/X5/M0_s
+ N_GND_X0/X2/M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13
mX31/X5/M1 N_VDD_X31/X5/M1_d N_X31/6_X31/X5/M1_g N_X31/5_X31/X5/M1_s
+ N_VDD_X31/X5/M1_b p L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12
*
.include "sipo_32.pex.netlist.SIPO_32.pxi"
*
.ends
*
*
