* SPICE NETLIST
***************************************

.SUBCKT v VDD IN OUT GND
** N=4 EP=4 IP=0 FDC=2
* PORT VDD VDD -8000 34000 METAL1
* PORT IN IN 17000 34000 METAL1
* PORT OUT OUT 17000 -20000 METAL1
* PORT GND GND 26000 34000 METAL1
M0 GND IN OUT GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=23000 $Y=1000 $D=1
M1 VDD IN OUT VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-11000 $Y=1000 $D=0
.ENDS
***************************************
.SUBCKT sipo VAL VALN VDD OUT IN GND CLK
** N=9 EP=7 IP=16 FDC=10
* PORT VAL VAL 172000 -97500 METAL1
* PORT VALN VALN 172000 -162000 METAL1
* PORT VDD VDD 205250 -240500 METAL1
* PORT VDD VDD 220750 110000 METAL1
* PORT OUT OUT 259500 -240000 METAL1
* PORT IN IN 259500 113000 METAL1
* PORT GND GND 283250 -241000 METAL1
* PORT GND GND 289250 113000 METAL1
* PORT CLK CLK 292000 52500 METAL1
* PORT CLK CLK 300000 -240000 METAL1
* PORT CLK CLK 315000 113000 METAL1
M0 IN CLK 6 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=265500 $Y=51500 $D=1
M1 IN CLK 6 VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=231500 $Y=51500 $D=0
X2 VDD VALN OUT GND v $T=242500 -199500 0 0 $X=222500 $Y=-221500
X3 VDD VAL VALN GND v $T=242500 -136000 0 0 $X=222500 $Y=-158000
X4 VDD 5 VAL GND v $T=242500 -74500 0 0 $X=222500 $Y=-96500
X5 VDD 6 5 GND v $T=242500 -12000 0 0 $X=222500 $Y=-34000
.ENDS
***************************************
.SUBCKT sipo_32 CLKN A3 A7 A11 A15 A19 A23 A27 A31 A0N A0 A1N A1 A2N A2 A3N A4N A4 A5N A5
+ A6N A6 A7N A8N A8 A9N A9 A10N A10 A11N A12N A12 A13N A13 A14N A14 A15N A16N A16 A17N
+ A17 A18N A18 A19N A20N A20 A21N A21 A22N A22 A23N A24N A24 A25N A25 A26N A26 A27N A28N A28
+ A29N A29 A30N A30 A31N VDD DIN GND CLK
** N=102 EP=69 IP=224 FDC=320
* PORT CLKN CLKN 380000 165000 METAL1
* PORT A3 A3 182000 -10311500 METAL1
* PORT A7 A7 182000 -8844000 METAL1
* PORT A11 A11 182000 -7384500 METAL1
* PORT A15 A15 182000 -5917000 METAL1
* PORT A19 A19 182000 -4458000 METAL1
* PORT A23 A23 182000 -2990500 METAL1
* PORT A27 A27 182000 -1531000 METAL1
* PORT A31 A31 182000 -63500 METAL1
* PORT A0N A0N 182500 -11474500 METAL1
* PORT A0 A0 182500 -11410000 METAL1
* PORT A1N A1N 182500 -11110000 METAL1
* PORT A1 A1 182500 -11045500 METAL1
* PORT A2N A2N 182500 -10740500 METAL1
* PORT A2 A2 182500 -10676000 METAL1
* PORT A3N A3N 182500 -10376000 METAL1
* PORT A4N A4N 182500 -10007000 METAL1
* PORT A4 A4 182500 -9942500 METAL1
* PORT A5N A5N 182500 -9642500 METAL1
* PORT A5 A5 182500 -9578000 METAL1
* PORT A6N A6N 182500 -9273000 METAL1
* PORT A6 A6 182500 -9208500 METAL1
* PORT A7N A7N 182500 -8908500 METAL1
* PORT A8N A8N 182500 -8547500 METAL1
* PORT A8 A8 182500 -8483000 METAL1
* PORT A9N A9N 182500 -8183000 METAL1
* PORT A9 A9 182500 -8118500 METAL1
* PORT A10N A10N 182500 -7813500 METAL1
* PORT A10 A10 182500 -7749000 METAL1
* PORT A11N A11N 182500 -7449000 METAL1
* PORT A12N A12N 182500 -7080000 METAL1
* PORT A12 A12 182500 -7015500 METAL1
* PORT A13N A13N 182500 -6715500 METAL1
* PORT A13 A13 182500 -6651000 METAL1
* PORT A14N A14N 182500 -6346000 METAL1
* PORT A14 A14 182500 -6281500 METAL1
* PORT A15N A15N 182500 -5981500 METAL1
* PORT A16N A16N 182500 -5621000 METAL1
* PORT A16 A16 182500 -5556500 METAL1
* PORT A17N A17N 182500 -5256500 METAL1
* PORT A17 A17 182500 -5192000 METAL1
* PORT A18N A18N 182500 -4887000 METAL1
* PORT A18 A18 182500 -4822500 METAL1
* PORT A19N A19N 182500 -4522500 METAL1
* PORT A20N A20N 182500 -4153500 METAL1
* PORT A20 A20 182500 -4089000 METAL1
* PORT A21N A21N 182500 -3789000 METAL1
* PORT A21 A21 182500 -3724500 METAL1
* PORT A22N A22N 182500 -3419500 METAL1
* PORT A22 A22 182500 -3355000 METAL1
* PORT A23N A23N 182500 -3055000 METAL1
* PORT A24N A24N 182500 -2694000 METAL1
* PORT A24 A24 182500 -2629500 METAL1
* PORT A25N A25N 182500 -2329500 METAL1
* PORT A25 A25 182500 -2265000 METAL1
* PORT A26N A26N 182500 -1960000 METAL1
* PORT A26 A26 182500 -1895500 METAL1
* PORT A27N A27N 182500 -1595500 METAL1
* PORT A28N A28N 182500 -1226500 METAL1
* PORT A28 A28 182500 -1162000 METAL1
* PORT A29N A29N 182500 -862000 METAL1
* PORT A29 A29 182500 -797500 METAL1
* PORT A30N A30N 182500 -492500 METAL1
* PORT A30 A30 182500 -428000 METAL1
* PORT A31N A31N 182500 -128000 METAL1
* PORT VDD VDD 245250 -11553000 METAL1
* PORT VDD VDD 260750 164750 METAL1
* PORT DIN DIN 299500 165000 METAL1
* PORT GND GND 323250 -11553500 METAL1
* PORT GND GND 329250 165250 METAL1
* PORT CLK CLK 355000 165000 METAL1
X0 A0 A0N VDD 102 68 GND CLKN sipo $T=40000 -11312500 0 0 $X=210000 $Y=-11554500
X1 A1 A1N VDD 68 69 GND CLK sipo $T=40000 -10948000 0 0 $X=210000 $Y=-11190000
X2 A2 A2N VDD 69 70 GND CLKN sipo $T=40000 -10578500 0 0 $X=210000 $Y=-10820500
X3 A3 A3N VDD 70 71 GND CLK sipo $T=40000 -10214000 0 0 $X=210000 $Y=-10456000
X4 A4 A4N VDD 71 72 GND CLKN sipo $T=40000 -9845000 0 0 $X=210000 $Y=-10087000
X5 A5 A5N VDD 72 73 GND CLK sipo $T=40000 -9480500 0 0 $X=210000 $Y=-9722500
X6 A6 A6N VDD 73 74 GND CLKN sipo $T=40000 -9111000 0 0 $X=210000 $Y=-9353000
X7 A7 A7N VDD 74 75 GND CLK sipo $T=40000 -8746500 0 0 $X=210000 $Y=-8988500
X8 A8 A8N VDD 75 76 GND CLKN sipo $T=40000 -8385500 0 0 $X=210000 $Y=-8627500
X9 A9 A9N VDD 76 77 GND CLK sipo $T=40000 -8021000 0 0 $X=210000 $Y=-8263000
X10 A10 A10N VDD 77 78 GND CLKN sipo $T=40000 -7651500 0 0 $X=210000 $Y=-7893500
X11 A11 A11N VDD 78 79 GND CLK sipo $T=40000 -7287000 0 0 $X=210000 $Y=-7529000
X12 A12 A12N VDD 79 80 GND CLKN sipo $T=40000 -6918000 0 0 $X=210000 $Y=-7160000
X13 A13 A13N VDD 80 81 GND CLK sipo $T=40000 -6553500 0 0 $X=210000 $Y=-6795500
X14 A14 A14N VDD 81 82 GND CLKN sipo $T=40000 -6184000 0 0 $X=210000 $Y=-6426000
X15 A15 A15N VDD 82 83 GND CLK sipo $T=40000 -5819500 0 0 $X=210000 $Y=-6061500
X16 A16 A16N VDD 83 84 GND CLKN sipo $T=40000 -5459000 0 0 $X=210000 $Y=-5701000
X17 A17 A17N VDD 84 85 GND CLK sipo $T=40000 -5094500 0 0 $X=210000 $Y=-5336500
X18 A18 A18N VDD 85 86 GND CLKN sipo $T=40000 -4725000 0 0 $X=210000 $Y=-4967000
X19 A19 A19N VDD 86 87 GND CLK sipo $T=40000 -4360500 0 0 $X=210000 $Y=-4602500
X20 A20 A20N VDD 87 88 GND CLKN sipo $T=40000 -3991500 0 0 $X=210000 $Y=-4233500
X21 A21 A21N VDD 88 89 GND CLK sipo $T=40000 -3627000 0 0 $X=210000 $Y=-3869000
X22 A22 A22N VDD 89 90 GND CLKN sipo $T=40000 -3257500 0 0 $X=210000 $Y=-3499500
X23 A23 A23N VDD 90 91 GND CLK sipo $T=40000 -2893000 0 0 $X=210000 $Y=-3135000
X24 A24 A24N VDD 91 92 GND CLKN sipo $T=40000 -2532000 0 0 $X=210000 $Y=-2774000
X25 A25 A25N VDD 92 93 GND CLK sipo $T=40000 -2167500 0 0 $X=210000 $Y=-2409500
X26 A26 A26N VDD 93 94 GND CLKN sipo $T=40000 -1798000 0 0 $X=210000 $Y=-2040000
X27 A27 A27N VDD 94 95 GND CLK sipo $T=40000 -1433500 0 0 $X=210000 $Y=-1675500
X28 A28 A28N VDD 95 96 GND CLKN sipo $T=40000 -1064500 0 0 $X=210000 $Y=-1306500
X29 A29 A29N VDD 96 97 GND CLK sipo $T=40000 -700000 0 0 $X=210000 $Y=-942000
X30 A30 A30N VDD 97 98 GND CLKN sipo $T=40000 -330500 0 0 $X=210000 $Y=-572500
X31 A31 A31N VDD 98 DIN GND CLK sipo $T=40000 34000 0 0 $X=210000 $Y=-208000
.ENDS
***************************************
