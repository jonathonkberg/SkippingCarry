* File: carry_skip_adder.pex.netlist
* Created: Sun Dec 18 19:16:29 2022
* Program "Calibre xRC"
* Version "v2012.2_36.25"
* 
.include /afs/cad/u/j/k/jk526/github/SkippingCarry/pre_sim/technologies/mosistsmc180_pex.sp
.include "carry_skip_adder.pex.netlist.pex"
.subckt CARRY_SKIP_ADDER  CINN A1N A3N A0N A2N VDD CIN GND SUM1 SUM3 SUM0 SUM2
+ B1N B3N B0N B2N A1 A3 A0 A2 COUTN COUT B1 B3 B0 B2
* 
* B2	B2
* B0	B0
* B3	B3
* B1	B1
* COUT	COUT
* COUTN	COUTN
* A2	A2
* A0	A0
* A3	A3
* A1	A1
* B2N	B2N
* B0N	B0N
* B3N	B3N
* B1N	B1N
* SUM2	SUM2
* SUM0	SUM0
* SUM3	SUM3
* SUM1	SUM1
* GND	GND
* CIN	CIN
* VDD	VDD
* A2N	A2N
* A0N	A0N
* A3N	A3N
* A1N	A1N
* CINN	CINN
M0 N_GND_M0_d N_27_M0_g N_SUM1_M0_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M1 N_GND_M1_d N_28_M1_g N_SUM3_M1_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M2 N_GND_M2_d N_29_M2_g N_SUM0_M2_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M3 N_GND_M3_d N_30_M3_g N_SUM2_M3_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M4 N_80_M4_d N_15_M4_g N_27_M4_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
M5 N_GND_M5_d N_18_M5_g N_80_M5_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
M6 N_81_M6_d N_A0N_M6_g N_GND_M6_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
M7 N_27_M7_d N_3_M7_g N_81_M7_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=4.374e-13
+ AS=5.832e-13
M8 N_82_M8_d N_19_M8_g N_28_M8_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=4.374e-13
M9 N_GND_M9_d N_20_M9_g N_82_M9_s N_GND_M0_b n L=1.8e-07 W=5.4e-07 AD=5.832e-13
+ AS=5.832e-13
M10 N_83_M10_d N_A2N_M10_g N_GND_M10_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M11 N_28_M11_d N_4_M11_g N_83_M11_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M12 N_84_M12_d N_14_M12_g N_29_M12_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M13 N_GND_M13_d N_21_M13_g N_84_M13_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M14 N_85_M14_d N_CIN_M14_g N_GND_M14_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M15 N_29_M15_d N_CINN_M15_g N_85_M15_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M16 N_86_M16_d N_16_M16_g N_30_M16_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M17 N_GND_M17_d N_22_M17_g N_86_M17_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M18 N_87_M18_d N_A1N_M18_g N_GND_M18_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M19 N_30_M19_d N_5_M19_g N_87_M19_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M20 N_GND_M20_d N_47_M20_g N_18_M20_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M21 N_GND_M21_d N_49_M21_g N_20_M21_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M22 N_GND_M22_d N_51_M22_g N_21_M22_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M23 N_GND_M23_d N_53_M23_g N_22_M23_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M24 N_GND_M24_d N_35_M24_g N_47_M24_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M25 N_88_M25_d N_36_M25_g N_GND_M25_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M26 N_47_M26_d N_B1N_M26_g N_88_M26_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M27 N_GND_M27_d N_38_M27_g N_49_M27_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M28 N_89_M28_d N_39_M28_g N_GND_M28_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M29 N_49_M29_d N_B3N_M29_g N_89_M29_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M30 N_GND_M30_d N_41_M30_g N_51_M30_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M31 N_90_M31_d N_42_M31_g N_GND_M31_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M32 N_51_M32_d N_B0N_M32_g N_90_M32_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M33 N_GND_M33_d N_44_M33_g N_53_M33_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M34 N_91_M34_d N_45_M34_g N_GND_M34_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M35 N_53_M35_d N_B2N_M35_g N_91_M35_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M36 N_GND_M36_d N_35_M36_g N_A1_M36_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M37 N_GND_M37_d N_38_M37_g N_A3_M37_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M38 N_GND_M38_d N_41_M38_g N_A0_M38_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M39 N_GND_M39_d N_44_M39_g N_A2_M39_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M40 N_35_M40_d N_36_M40_g N_GND_M40_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M41 N_GND_M41_d N_B1N_M41_g N_35_M41_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M42 N_38_M42_d N_39_M42_g N_GND_M42_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M43 N_GND_M43_d N_B3N_M43_g N_38_M43_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M44 N_41_M44_d N_42_M44_g N_GND_M44_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M45 N_GND_M45_d N_B0N_M45_g N_41_M45_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M46 N_44_M46_d N_45_M46_g N_GND_M46_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M47 N_GND_M47_d N_B2N_M47_g N_44_M47_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M48 N_GND_M48_d N_5_M48_g N_A1N_M48_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M49 N_GND_M49_d N_2_M49_g N_A3N_M49_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M50 N_GND_M50_d N_3_M50_g N_A0N_M50_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M51 N_GND_M51_d N_4_M51_g N_A2N_M51_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M52 N_GND_M52_d N_COUTN_M52_g N_COUT_M52_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M53 N_92_M53_d N_36_M53_g N_5_M53_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M54 N_GND_M54_d N_B1N_M54_g N_92_M54_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M55 N_93_M55_d N_A1_M55_g N_GND_M55_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M56 N_5_M56_d N_A0N_M56_g N_93_M56_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M57 N_94_M57_d N_39_M57_g N_2_M57_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M58 N_GND_M58_d N_B3N_M58_g N_94_M58_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M59 N_95_M59_d N_A3_M59_g N_GND_M59_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M60 N_2_M60_d N_A2N_M60_g N_95_M60_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M61 N_96_M61_d N_42_M61_g N_3_M61_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M62 N_GND_M62_d N_B0N_M62_g N_96_M62_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M63 N_97_M63_d N_A0_M63_g N_GND_M63_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M64 N_3_M64_d N_CIN_M64_g N_97_M64_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M65 N_98_M65_d N_45_M65_g N_4_M65_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M66 N_GND_M66_d N_B2N_M66_g N_98_M66_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M67 N_99_M67_d N_A2_M67_g N_GND_M67_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M68 N_4_M68_d N_A1N_M68_g N_99_M68_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M69 N_100_M69_d N_59_M69_g N_COUTN_M69_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M70 N_GND_M70_d N_CIN_M70_g N_100_M70_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M71 N_101_M71_d N_A3N_M71_g N_GND_M71_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M72 N_COUTN_M72_d N_60_M72_g N_101_M72_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M73 N_GND_M73_d N_60_M73_g N_A3N_M73_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M74 N_102_M74_d N_14_M74_g N_GND_M74_s N_GND_M0_b n L=1.8e-07 W=2.16e-06
+ AD=2.3328e-12 AS=1.7496e-12
M75 N_103_M75_d N_15_M75_g N_102_M75_s N_GND_M0_b n L=1.8e-07 W=2.16e-06
+ AD=2.3328e-12 AS=2.3328e-12
M76 N_104_M76_d N_16_M76_g N_103_M76_s N_GND_M0_b n L=1.8e-07 W=2.16e-06
+ AD=2.3328e-12 AS=2.3328e-12
M77 N_60_M77_d N_19_M77_g N_104_M77_s N_GND_M0_b n L=1.8e-07 W=2.16e-06
+ AD=1.7496e-12 AS=2.3328e-12
M78 N_GND_M78_d N_76_M78_g N_15_M78_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M79 N_GND_M79_d N_77_M79_g N_19_M79_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M80 N_GND_M80_d N_78_M80_g N_14_M80_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M81 N_GND_M81_d N_79_M81_g N_16_M81_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=4.374e-13
M82 N_105_M82_d N_B1N_M82_g N_76_M82_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M83 N_GND_M83_d N_B1_M83_g N_105_M83_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M84 N_106_M84_d N_A1N_M84_g N_GND_M84_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M85 N_76_M85_d N_A1_M85_g N_106_M85_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M86 N_107_M86_d N_B3N_M86_g N_77_M86_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M87 N_GND_M87_d N_B3_M87_g N_107_M87_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M88 N_108_M88_d N_A3N_M88_g N_GND_M88_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M89 N_77_M89_d N_A3_M89_g N_108_M89_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M90 N_109_M90_d N_B0N_M90_g N_78_M90_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M91 N_GND_M91_d N_B0_M91_g N_109_M91_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M92 N_110_M92_d N_A0N_M92_g N_GND_M92_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M93 N_78_M93_d N_A0_M93_g N_110_M93_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M94 N_111_M94_d N_B2N_M94_g N_79_M94_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=4.374e-13
M95 N_GND_M95_d N_B2_M95_g N_111_M95_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M96 N_112_M96_d N_A2N_M96_g N_GND_M96_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=5.832e-13 AS=5.832e-13
M97 N_79_M97_d N_A2_M97_g N_112_M97_s N_GND_M0_b n L=1.8e-07 W=5.4e-07
+ AD=4.374e-13 AS=5.832e-13
M98 N_23_M98_d N_A0N_M98_g N_VDD_M98_s N_VDD_M98_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M99 N_27_M99_d N_15_M99_g N_23_M99_s N_VDD_M98_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M100 N_23_M100_d N_18_M100_g N_27_M100_s N_VDD_M98_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M101 N_VDD_M101_d N_3_M101_g N_23_M101_s N_VDD_M98_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M102 N_24_M102_d N_A2N_M102_g N_VDD_M102_s N_VDD_M102_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M103 N_28_M103_d N_19_M103_g N_24_M103_s N_VDD_M102_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M104 N_24_M104_d N_20_M104_g N_28_M104_s N_VDD_M102_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M105 N_VDD_M105_d N_4_M105_g N_24_M105_s N_VDD_M102_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M106 N_25_M106_d N_CIN_M106_g N_VDD_M106_s N_VDD_M106_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M107 N_29_M107_d N_14_M107_g N_25_M107_s N_VDD_M106_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M108 N_25_M108_d N_21_M108_g N_29_M108_s N_VDD_M106_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M109 N_VDD_M109_d N_CINN_M109_g N_25_M109_s N_VDD_M106_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M110 N_26_M110_d N_A1N_M110_g N_VDD_M110_s N_VDD_M110_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M111 N_30_M111_d N_16_M111_g N_26_M111_s N_VDD_M110_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M112 N_26_M112_d N_22_M112_g N_30_M112_s N_VDD_M110_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M113 N_VDD_M113_d N_5_M113_g N_26_M113_s N_VDD_M110_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M114 N_VDD_M114_d N_27_M114_g N_SUM1_M114_s N_VDD_M98_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M115 N_VDD_M115_d N_28_M115_g N_SUM3_M115_s N_VDD_M102_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M116 N_VDD_M116_d N_29_M116_g N_SUM0_M116_s N_VDD_M106_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M117 N_VDD_M117_d N_30_M117_g N_SUM2_M117_s N_VDD_M110_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M118 N_48_M118_d N_35_M118_g N_47_M118_s N_VDD_M118_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M119 N_VDD_M119_d N_36_M119_g N_48_M119_s N_VDD_M118_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M120 N_48_M120_d N_B1N_M120_g N_VDD_M120_s N_VDD_M118_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M121 N_50_M121_d N_38_M121_g N_49_M121_s N_VDD_M121_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M122 N_VDD_M122_d N_39_M122_g N_50_M122_s N_VDD_M121_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M123 N_50_M123_d N_B3N_M123_g N_VDD_M123_s N_VDD_M121_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M124 N_52_M124_d N_41_M124_g N_51_M124_s N_VDD_M124_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M125 N_VDD_M125_d N_42_M125_g N_52_M125_s N_VDD_M124_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M126 N_52_M126_d N_B0N_M126_g N_VDD_M126_s N_VDD_M124_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M127 N_54_M127_d N_44_M127_g N_53_M127_s N_VDD_M127_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M128 N_VDD_M128_d N_45_M128_g N_54_M128_s N_VDD_M127_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M129 N_54_M129_d N_B2N_M129_g N_VDD_M129_s N_VDD_M127_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M130 N_VDD_M130_d N_47_M130_g N_18_M130_s N_VDD_M118_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M131 N_VDD_M131_d N_49_M131_g N_20_M131_s N_VDD_M121_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M132 N_VDD_M132_d N_51_M132_g N_21_M132_s N_VDD_M124_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M133 N_VDD_M133_d N_53_M133_g N_22_M133_s N_VDD_M127_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M134 N_113_M134_d N_36_M134_g N_VDD_M134_s N_VDD_M134_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M135 N_35_M135_d N_B1N_M135_g N_113_M135_s N_VDD_M134_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M136 N_114_M136_d N_39_M136_g N_VDD_M136_s N_VDD_M136_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M137 N_38_M137_d N_B3N_M137_g N_114_M137_s N_VDD_M136_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M138 N_115_M138_d N_42_M138_g N_VDD_M138_s N_VDD_M138_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M139 N_41_M139_d N_B0N_M139_g N_115_M139_s N_VDD_M138_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M140 N_116_M140_d N_45_M140_g N_VDD_M140_s N_VDD_M140_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M141 N_44_M141_d N_B2N_M141_g N_116_M141_s N_VDD_M140_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M142 N_VDD_M142_d N_35_M142_g N_A1_M142_s N_VDD_M134_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M143 N_VDD_M143_d N_38_M143_g N_A3_M143_s N_VDD_M136_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M144 N_VDD_M144_d N_41_M144_g N_A0_M144_s N_VDD_M138_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M145 N_VDD_M145_d N_44_M145_g N_A2_M145_s N_VDD_M140_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M146 N_61_M146_d N_A1_M146_g N_VDD_M146_s N_VDD_M146_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M147 N_5_M147_d N_36_M147_g N_61_M147_s N_VDD_M146_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M148 N_61_M148_d N_B1N_M148_g N_5_M148_s N_VDD_M146_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M149 N_VDD_M149_d N_A0N_M149_g N_61_M149_s N_VDD_M146_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M150 N_62_M150_d N_A3_M150_g N_VDD_M150_s N_VDD_M150_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M151 N_2_M151_d N_39_M151_g N_62_M151_s N_VDD_M150_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M152 N_62_M152_d N_B3N_M152_g N_2_M152_s N_VDD_M150_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M153 N_VDD_M153_d N_A2N_M153_g N_62_M153_s N_VDD_M150_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M154 N_63_M154_d N_A0_M154_g N_VDD_M154_s N_VDD_M154_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M155 N_3_M155_d N_42_M155_g N_63_M155_s N_VDD_M154_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M156 N_63_M156_d N_B0N_M156_g N_3_M156_s N_VDD_M154_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M157 N_VDD_M157_d N_CIN_M157_g N_63_M157_s N_VDD_M154_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M158 N_64_M158_d N_A2_M158_g N_VDD_M158_s N_VDD_M158_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M159 N_4_M159_d N_45_M159_g N_64_M159_s N_VDD_M158_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M160 N_64_M160_d N_B2N_M160_g N_4_M160_s N_VDD_M158_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M161 N_VDD_M161_d N_A1N_M161_g N_64_M161_s N_VDD_M158_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M162 N_65_M162_d N_A3N_M162_g N_11_M162_s N_11_M162_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M163 N_COUTN_M163_d N_59_M163_g N_65_M163_s N_11_M162_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M164 N_65_M164_d N_CIN_M164_g N_COUTN_M164_s N_11_M162_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M165 N_11_M165_d N_60_M165_g N_65_M165_s N_11_M162_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M166 N_VDD_M166_d N_5_M166_g N_A1N_M166_s N_VDD_M146_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M167 N_VDD_M167_d N_2_M167_g N_A3N_M167_s N_VDD_M150_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M168 N_VDD_M168_d N_3_M168_g N_A0N_M168_s N_VDD_M154_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M169 N_VDD_M169_d N_4_M169_g N_A2N_M169_s N_VDD_M158_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M170 N_11_M170_d N_COUTN_M170_g N_COUT_M170_s N_11_M162_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M171 N_72_M171_d N_A1N_M171_g N_VDD_M171_s N_VDD_M171_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M172 N_76_M172_d N_B1N_M172_g N_72_M172_s N_VDD_M171_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M173 N_72_M173_d N_B1_M173_g N_76_M173_s N_VDD_M171_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M174 N_VDD_M174_d N_A1_M174_g N_72_M174_s N_VDD_M171_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M175 N_73_M175_d N_A3N_M175_g N_VDD_M175_s N_VDD_M175_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M176 N_77_M176_d N_B3N_M176_g N_73_M176_s N_VDD_M175_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M177 N_73_M177_d N_B3_M177_g N_77_M177_s N_VDD_M175_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M178 N_VDD_M178_d N_A3_M178_g N_73_M178_s N_VDD_M175_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M179 N_74_M179_d N_A0N_M179_g N_VDD_M179_s N_VDD_M179_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M180 N_78_M180_d N_B0N_M180_g N_74_M180_s N_VDD_M179_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M181 N_74_M181_d N_B0_M181_g N_78_M181_s N_VDD_M179_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M182 N_VDD_M182_d N_A0_M182_g N_74_M182_s N_VDD_M179_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M183 N_75_M183_d N_A2N_M183_g N_VDD_M183_s N_VDD_M183_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=2.3328e-12
M184 N_79_M184_d N_B2N_M184_g N_75_M184_s N_VDD_M183_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M185 N_75_M185_d N_B2_M185_g N_79_M185_s N_VDD_M183_b p L=1.8e-07 W=2.88e-06
+ AD=3.1104e-12 AS=3.1104e-12
M186 N_VDD_M186_d N_A2_M186_g N_75_M186_s N_VDD_M183_b p L=1.8e-07 W=2.88e-06
+ AD=2.3328e-12 AS=3.1104e-12
M187 N_13_M187_d N_60_M187_g N_A3N_M187_s N_13_M187_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M188 N_60_M188_d N_14_M188_g N_13_M188_s N_13_M187_b p L=1.8e-07 W=1.44e-06
+ AD=1.5552e-12 AS=1.1664e-12
M189 N_13_M189_d N_15_M189_g N_60_M189_s N_13_M187_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.5552e-12
M190 N_60_M190_d N_16_M190_g N_13_M190_s N_13_M187_b p L=1.8e-07 W=1.44e-06
+ AD=1.5552e-12 AS=1.1664e-12
M191 N_13_M191_d N_19_M191_g N_60_M191_s N_13_M187_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.5552e-12
M192 N_VDD_M192_d N_76_M192_g N_15_M192_s N_VDD_M171_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M193 N_VDD_M193_d N_77_M193_g N_19_M193_s N_VDD_M175_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M194 N_VDD_M194_d N_78_M194_g N_14_M194_s N_VDD_M179_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
M195 N_VDD_M195_d N_79_M195_g N_16_M195_s N_VDD_M183_b p L=1.8e-07 W=1.44e-06
+ AD=1.1664e-12 AS=1.1664e-12
*
.include "carry_skip_adder.pex.netlist.CARRY_SKIP_ADDER.pxi"
*
.ends
*
*
