* SPICE NETLIST
***************************************

.SUBCKT three_in_aoi VDD Y C B A GND
** N=8 EP=6 IP=0 FDC=6
* PORT VDD VDD -20000 37000 METAL1
* PORT Y Y 50000 -8000 METAL1
* PORT C C 73000 -1000 METAL1
* PORT B B 89000 30000 METAL1
* PORT A A 89000 44000 METAL1
* PORT GND GND 86000 3000 METAL1
M0 GND C Y GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=4.374e-13 $X=62000 $Y=15000 $D=1
M1 8 B GND GND N L=1.8e-07 W=5.4e-07 AD=5.832e-13 AS=5.832e-13 $X=62000 $Y=29000 $D=1
M2 Y A 8 GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=5.832e-13 $X=62000 $Y=43000 $D=1
M3 2 C Y VDD P L=1.8e-07 W=1.53e-06 AD=1.6524e-12 AS=1.2393e-12 $X=18000 $Y=15000 $D=0
M4 VDD B 2 VDD P L=1.8e-07 W=1.53e-06 AD=1.6524e-12 AS=1.6524e-12 $X=18000 $Y=29000 $D=0
M5 2 A VDD VDD P L=1.8e-07 W=1.53e-06 AD=1.2393e-12 AS=1.6524e-12 $X=18000 $Y=43000 $D=0
.ENDS
***************************************
