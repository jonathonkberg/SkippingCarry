* SPICE NETLIST
***************************************

.SUBCKT base_inverter VDD IN OUT GND
** N=4 EP=4 IP=0 FDC=2
* PORT VDD VDD 1000 44000 METAL1
* PORT IN IN 26000 44000 METAL1
* PORT OUT OUT 26000 -10000 METAL1
* PORT GND GND 35000 44000 METAL1
M0 GND IN OUT GND N L=1.8e-07 W=5.4e-07 AD=4.374e-13 AS=4.374e-13 $X=32000 $Y=11000 $D=1
M1 VDD IN OUT VDD P L=1.8e-07 W=1.44e-06 AD=1.1664e-12 AS=1.1664e-12 $X=-2000 $Y=11000 $D=0
.ENDS
***************************************
